
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h45e8c2b2;
    ram_cell[       1] = 32'h0;  // 32'ha0e37c50;
    ram_cell[       2] = 32'h0;  // 32'h40a42c52;
    ram_cell[       3] = 32'h0;  // 32'h0cbb4e15;
    ram_cell[       4] = 32'h0;  // 32'hf6cc8129;
    ram_cell[       5] = 32'h0;  // 32'hfe7b3942;
    ram_cell[       6] = 32'h0;  // 32'h24eccbc3;
    ram_cell[       7] = 32'h0;  // 32'h268dd8ee;
    ram_cell[       8] = 32'h0;  // 32'h8d215f19;
    ram_cell[       9] = 32'h0;  // 32'h87485cd6;
    ram_cell[      10] = 32'h0;  // 32'h39bc467b;
    ram_cell[      11] = 32'h0;  // 32'h7bdc805d;
    ram_cell[      12] = 32'h0;  // 32'h97a50d6c;
    ram_cell[      13] = 32'h0;  // 32'h458936bc;
    ram_cell[      14] = 32'h0;  // 32'h8b7fa195;
    ram_cell[      15] = 32'h0;  // 32'h7ab2f074;
    ram_cell[      16] = 32'h0;  // 32'h124e7d8a;
    ram_cell[      17] = 32'h0;  // 32'hf9756787;
    ram_cell[      18] = 32'h0;  // 32'hd3e65800;
    ram_cell[      19] = 32'h0;  // 32'h559bc980;
    ram_cell[      20] = 32'h0;  // 32'h52468ded;
    ram_cell[      21] = 32'h0;  // 32'h0ac2461d;
    ram_cell[      22] = 32'h0;  // 32'h9d59c195;
    ram_cell[      23] = 32'h0;  // 32'h4bfd277f;
    ram_cell[      24] = 32'h0;  // 32'hf4c05c82;
    ram_cell[      25] = 32'h0;  // 32'h3db632f6;
    ram_cell[      26] = 32'h0;  // 32'h019c2cdb;
    ram_cell[      27] = 32'h0;  // 32'h457f70a0;
    ram_cell[      28] = 32'h0;  // 32'h1c191151;
    ram_cell[      29] = 32'h0;  // 32'h5bb71630;
    ram_cell[      30] = 32'h0;  // 32'h827bd456;
    ram_cell[      31] = 32'h0;  // 32'h1fb5fadd;
    ram_cell[      32] = 32'h0;  // 32'h6dd5e0b2;
    ram_cell[      33] = 32'h0;  // 32'hf623916a;
    ram_cell[      34] = 32'h0;  // 32'h2e9ddced;
    ram_cell[      35] = 32'h0;  // 32'h1baed27f;
    ram_cell[      36] = 32'h0;  // 32'h64f0042f;
    ram_cell[      37] = 32'h0;  // 32'h4a55f4e1;
    ram_cell[      38] = 32'h0;  // 32'hb7d0ccab;
    ram_cell[      39] = 32'h0;  // 32'heabea5cf;
    ram_cell[      40] = 32'h0;  // 32'hd83772f8;
    ram_cell[      41] = 32'h0;  // 32'h18133ff3;
    ram_cell[      42] = 32'h0;  // 32'h4c8ae3c7;
    ram_cell[      43] = 32'h0;  // 32'hcb7b7ef6;
    ram_cell[      44] = 32'h0;  // 32'he6689cc3;
    ram_cell[      45] = 32'h0;  // 32'h1bd42672;
    ram_cell[      46] = 32'h0;  // 32'hff464453;
    ram_cell[      47] = 32'h0;  // 32'hd8599bd2;
    ram_cell[      48] = 32'h0;  // 32'h96aed738;
    ram_cell[      49] = 32'h0;  // 32'h99f63909;
    ram_cell[      50] = 32'h0;  // 32'hdfeeb6ce;
    ram_cell[      51] = 32'h0;  // 32'he74a50d5;
    ram_cell[      52] = 32'h0;  // 32'ha4845fe0;
    ram_cell[      53] = 32'h0;  // 32'h18cdba80;
    ram_cell[      54] = 32'h0;  // 32'hda3a8543;
    ram_cell[      55] = 32'h0;  // 32'h5e1eed87;
    ram_cell[      56] = 32'h0;  // 32'h18cf43a1;
    ram_cell[      57] = 32'h0;  // 32'h7e1aa9cf;
    ram_cell[      58] = 32'h0;  // 32'h3604fb89;
    ram_cell[      59] = 32'h0;  // 32'hb54fd431;
    ram_cell[      60] = 32'h0;  // 32'he2cef799;
    ram_cell[      61] = 32'h0;  // 32'had150635;
    ram_cell[      62] = 32'h0;  // 32'hb21feb7a;
    ram_cell[      63] = 32'h0;  // 32'h4d816d37;
    ram_cell[      64] = 32'h0;  // 32'he1b63d0f;
    ram_cell[      65] = 32'h0;  // 32'h3448dc1f;
    ram_cell[      66] = 32'h0;  // 32'h86a60d7b;
    ram_cell[      67] = 32'h0;  // 32'hc573a294;
    ram_cell[      68] = 32'h0;  // 32'hff21539c;
    ram_cell[      69] = 32'h0;  // 32'h419f472e;
    ram_cell[      70] = 32'h0;  // 32'h40faec76;
    ram_cell[      71] = 32'h0;  // 32'h62e4c8c7;
    ram_cell[      72] = 32'h0;  // 32'h65c41fa7;
    ram_cell[      73] = 32'h0;  // 32'h9e9fe45f;
    ram_cell[      74] = 32'h0;  // 32'h8f9a3be0;
    ram_cell[      75] = 32'h0;  // 32'he2a3c28f;
    ram_cell[      76] = 32'h0;  // 32'h3f6a651e;
    ram_cell[      77] = 32'h0;  // 32'h12d25cc8;
    ram_cell[      78] = 32'h0;  // 32'h87216a79;
    ram_cell[      79] = 32'h0;  // 32'h0cfdc85f;
    ram_cell[      80] = 32'h0;  // 32'hd4623dc9;
    ram_cell[      81] = 32'h0;  // 32'h339f7d75;
    ram_cell[      82] = 32'h0;  // 32'h0cd89e54;
    ram_cell[      83] = 32'h0;  // 32'h8cb80d2e;
    ram_cell[      84] = 32'h0;  // 32'h15870643;
    ram_cell[      85] = 32'h0;  // 32'h66a9626c;
    ram_cell[      86] = 32'h0;  // 32'h4fd6012f;
    ram_cell[      87] = 32'h0;  // 32'h0841d17e;
    ram_cell[      88] = 32'h0;  // 32'h5c2415fa;
    ram_cell[      89] = 32'h0;  // 32'h628272e7;
    ram_cell[      90] = 32'h0;  // 32'ha8a57310;
    ram_cell[      91] = 32'h0;  // 32'hdc943185;
    ram_cell[      92] = 32'h0;  // 32'h834372cb;
    ram_cell[      93] = 32'h0;  // 32'he4c9ffe2;
    ram_cell[      94] = 32'h0;  // 32'h48270933;
    ram_cell[      95] = 32'h0;  // 32'hd94eb740;
    ram_cell[      96] = 32'h0;  // 32'hde596e15;
    ram_cell[      97] = 32'h0;  // 32'h5f34d0d6;
    ram_cell[      98] = 32'h0;  // 32'h288fe1c3;
    ram_cell[      99] = 32'h0;  // 32'hdda2a235;
    ram_cell[     100] = 32'h0;  // 32'h0a91fa21;
    ram_cell[     101] = 32'h0;  // 32'h02958ff0;
    ram_cell[     102] = 32'h0;  // 32'h63b81525;
    ram_cell[     103] = 32'h0;  // 32'h581886c6;
    ram_cell[     104] = 32'h0;  // 32'h035e2d7d;
    ram_cell[     105] = 32'h0;  // 32'ha29d5e79;
    ram_cell[     106] = 32'h0;  // 32'h644418f6;
    ram_cell[     107] = 32'h0;  // 32'hb2380809;
    ram_cell[     108] = 32'h0;  // 32'h9d2f1687;
    ram_cell[     109] = 32'h0;  // 32'h8cccb089;
    ram_cell[     110] = 32'h0;  // 32'h52783f05;
    ram_cell[     111] = 32'h0;  // 32'hfe15eaab;
    ram_cell[     112] = 32'h0;  // 32'h13dda05a;
    ram_cell[     113] = 32'h0;  // 32'h2c9a3a83;
    ram_cell[     114] = 32'h0;  // 32'hb2a963c4;
    ram_cell[     115] = 32'h0;  // 32'hadf5b875;
    ram_cell[     116] = 32'h0;  // 32'h09447dca;
    ram_cell[     117] = 32'h0;  // 32'hcb80071f;
    ram_cell[     118] = 32'h0;  // 32'hc2320cf0;
    ram_cell[     119] = 32'h0;  // 32'h67c97b61;
    ram_cell[     120] = 32'h0;  // 32'hbd23139f;
    ram_cell[     121] = 32'h0;  // 32'hc467cf88;
    ram_cell[     122] = 32'h0;  // 32'h3844d396;
    ram_cell[     123] = 32'h0;  // 32'hedf3d39a;
    ram_cell[     124] = 32'h0;  // 32'h2952bd4e;
    ram_cell[     125] = 32'h0;  // 32'h549d917e;
    ram_cell[     126] = 32'h0;  // 32'h07872ad4;
    ram_cell[     127] = 32'h0;  // 32'h1864ea4b;
    ram_cell[     128] = 32'h0;  // 32'h56bc5ced;
    ram_cell[     129] = 32'h0;  // 32'h4b0a8a6d;
    ram_cell[     130] = 32'h0;  // 32'he37ee270;
    ram_cell[     131] = 32'h0;  // 32'he211489b;
    ram_cell[     132] = 32'h0;  // 32'hbb1b2ec8;
    ram_cell[     133] = 32'h0;  // 32'h24cab396;
    ram_cell[     134] = 32'h0;  // 32'hd5129929;
    ram_cell[     135] = 32'h0;  // 32'h92355c68;
    ram_cell[     136] = 32'h0;  // 32'hddedf773;
    ram_cell[     137] = 32'h0;  // 32'h94ea136a;
    ram_cell[     138] = 32'h0;  // 32'h91e5e47f;
    ram_cell[     139] = 32'h0;  // 32'hfe6c051e;
    ram_cell[     140] = 32'h0;  // 32'h54bb090a;
    ram_cell[     141] = 32'h0;  // 32'hc589cacc;
    ram_cell[     142] = 32'h0;  // 32'hab50c00c;
    ram_cell[     143] = 32'h0;  // 32'hf1a09bf1;
    ram_cell[     144] = 32'h0;  // 32'hde7e9dd0;
    ram_cell[     145] = 32'h0;  // 32'h0351885c;
    ram_cell[     146] = 32'h0;  // 32'h95ef0b6c;
    ram_cell[     147] = 32'h0;  // 32'h10710574;
    ram_cell[     148] = 32'h0;  // 32'h7bda552e;
    ram_cell[     149] = 32'h0;  // 32'h8fb9ce0e;
    ram_cell[     150] = 32'h0;  // 32'hd323db3e;
    ram_cell[     151] = 32'h0;  // 32'h1a9f4e3e;
    ram_cell[     152] = 32'h0;  // 32'h1c400503;
    ram_cell[     153] = 32'h0;  // 32'h4b2f63cb;
    ram_cell[     154] = 32'h0;  // 32'hdb93e493;
    ram_cell[     155] = 32'h0;  // 32'hc87f34dc;
    ram_cell[     156] = 32'h0;  // 32'hd7ea49cf;
    ram_cell[     157] = 32'h0;  // 32'h5d3637b8;
    ram_cell[     158] = 32'h0;  // 32'h3e44fd52;
    ram_cell[     159] = 32'h0;  // 32'heb443a30;
    ram_cell[     160] = 32'h0;  // 32'h9deb9457;
    ram_cell[     161] = 32'h0;  // 32'h76212144;
    ram_cell[     162] = 32'h0;  // 32'h29b3d15a;
    ram_cell[     163] = 32'h0;  // 32'h90293e2e;
    ram_cell[     164] = 32'h0;  // 32'h29e3cd84;
    ram_cell[     165] = 32'h0;  // 32'h45c88b1b;
    ram_cell[     166] = 32'h0;  // 32'hc957f916;
    ram_cell[     167] = 32'h0;  // 32'hfdce0116;
    ram_cell[     168] = 32'h0;  // 32'h83be1a03;
    ram_cell[     169] = 32'h0;  // 32'h05438023;
    ram_cell[     170] = 32'h0;  // 32'h7722550f;
    ram_cell[     171] = 32'h0;  // 32'h0835b060;
    ram_cell[     172] = 32'h0;  // 32'h2dd68581;
    ram_cell[     173] = 32'h0;  // 32'hef3f0b72;
    ram_cell[     174] = 32'h0;  // 32'he80694c6;
    ram_cell[     175] = 32'h0;  // 32'h4a841642;
    ram_cell[     176] = 32'h0;  // 32'hc2728213;
    ram_cell[     177] = 32'h0;  // 32'h186bb0f0;
    ram_cell[     178] = 32'h0;  // 32'hb2c9e570;
    ram_cell[     179] = 32'h0;  // 32'haa77884b;
    ram_cell[     180] = 32'h0;  // 32'h941e0f34;
    ram_cell[     181] = 32'h0;  // 32'h8d7a9ef3;
    ram_cell[     182] = 32'h0;  // 32'he8ecd89d;
    ram_cell[     183] = 32'h0;  // 32'hd6dfa0f8;
    ram_cell[     184] = 32'h0;  // 32'h3a8fe9eb;
    ram_cell[     185] = 32'h0;  // 32'h6428bf55;
    ram_cell[     186] = 32'h0;  // 32'hde99d5d7;
    ram_cell[     187] = 32'h0;  // 32'h3b7462fa;
    ram_cell[     188] = 32'h0;  // 32'he835fbbb;
    ram_cell[     189] = 32'h0;  // 32'hc9a71fb5;
    ram_cell[     190] = 32'h0;  // 32'h3d054c6b;
    ram_cell[     191] = 32'h0;  // 32'hd7d0687f;
    ram_cell[     192] = 32'h0;  // 32'ha84cdb0d;
    ram_cell[     193] = 32'h0;  // 32'heb26249b;
    ram_cell[     194] = 32'h0;  // 32'he1f5d733;
    ram_cell[     195] = 32'h0;  // 32'hfb0ed7fd;
    ram_cell[     196] = 32'h0;  // 32'h87cc5eb1;
    ram_cell[     197] = 32'h0;  // 32'h5d3d46bd;
    ram_cell[     198] = 32'h0;  // 32'he09290f4;
    ram_cell[     199] = 32'h0;  // 32'hbeb4efc6;
    ram_cell[     200] = 32'h0;  // 32'h31be8edd;
    ram_cell[     201] = 32'h0;  // 32'h47362498;
    ram_cell[     202] = 32'h0;  // 32'he170639f;
    ram_cell[     203] = 32'h0;  // 32'hdeb41c2a;
    ram_cell[     204] = 32'h0;  // 32'h9b59885b;
    ram_cell[     205] = 32'h0;  // 32'hcff4075c;
    ram_cell[     206] = 32'h0;  // 32'ha2eb6c2c;
    ram_cell[     207] = 32'h0;  // 32'hc2e33e17;
    ram_cell[     208] = 32'h0;  // 32'he6187482;
    ram_cell[     209] = 32'h0;  // 32'ha50cb1ec;
    ram_cell[     210] = 32'h0;  // 32'h899aad95;
    ram_cell[     211] = 32'h0;  // 32'h7bfa24af;
    ram_cell[     212] = 32'h0;  // 32'h086249af;
    ram_cell[     213] = 32'h0;  // 32'h64dbdf88;
    ram_cell[     214] = 32'h0;  // 32'h4eefca52;
    ram_cell[     215] = 32'h0;  // 32'h7503a2d4;
    ram_cell[     216] = 32'h0;  // 32'h21c2c978;
    ram_cell[     217] = 32'h0;  // 32'h76734d0e;
    ram_cell[     218] = 32'h0;  // 32'ha67c4a61;
    ram_cell[     219] = 32'h0;  // 32'h1ef71313;
    ram_cell[     220] = 32'h0;  // 32'h1c5ee2f3;
    ram_cell[     221] = 32'h0;  // 32'h2f4c2b66;
    ram_cell[     222] = 32'h0;  // 32'ha53fc993;
    ram_cell[     223] = 32'h0;  // 32'h62604652;
    ram_cell[     224] = 32'h0;  // 32'hf39a83cd;
    ram_cell[     225] = 32'h0;  // 32'h4c3685fb;
    ram_cell[     226] = 32'h0;  // 32'ha42ee5ee;
    ram_cell[     227] = 32'h0;  // 32'h5943b230;
    ram_cell[     228] = 32'h0;  // 32'hf9a8569b;
    ram_cell[     229] = 32'h0;  // 32'h58dc8408;
    ram_cell[     230] = 32'h0;  // 32'h347ac094;
    ram_cell[     231] = 32'h0;  // 32'hcc4b7145;
    ram_cell[     232] = 32'h0;  // 32'had5fce0d;
    ram_cell[     233] = 32'h0;  // 32'h8345bbc9;
    ram_cell[     234] = 32'h0;  // 32'h85b9e208;
    ram_cell[     235] = 32'h0;  // 32'h11525b49;
    ram_cell[     236] = 32'h0;  // 32'heecdbd2e;
    ram_cell[     237] = 32'h0;  // 32'hf36ee2d5;
    ram_cell[     238] = 32'h0;  // 32'h74f2ce44;
    ram_cell[     239] = 32'h0;  // 32'haed0a135;
    ram_cell[     240] = 32'h0;  // 32'h01469a6c;
    ram_cell[     241] = 32'h0;  // 32'hbba6bc21;
    ram_cell[     242] = 32'h0;  // 32'h096611f2;
    ram_cell[     243] = 32'h0;  // 32'hc1fea6e5;
    ram_cell[     244] = 32'h0;  // 32'h1f8fa7e4;
    ram_cell[     245] = 32'h0;  // 32'hf8c900a6;
    ram_cell[     246] = 32'h0;  // 32'h24b2395e;
    ram_cell[     247] = 32'h0;  // 32'h437f70e8;
    ram_cell[     248] = 32'h0;  // 32'hc70e8a46;
    ram_cell[     249] = 32'h0;  // 32'he951d811;
    ram_cell[     250] = 32'h0;  // 32'h36834189;
    ram_cell[     251] = 32'h0;  // 32'h4103e2ba;
    ram_cell[     252] = 32'h0;  // 32'hd50de9f2;
    ram_cell[     253] = 32'h0;  // 32'hb9230823;
    ram_cell[     254] = 32'h0;  // 32'he512cc29;
    ram_cell[     255] = 32'h0;  // 32'hed699b28;
    ram_cell[     256] = 32'h0;  // 32'hfa24d840;
    ram_cell[     257] = 32'h0;  // 32'he354bf8d;
    ram_cell[     258] = 32'h0;  // 32'h5a48a849;
    ram_cell[     259] = 32'h0;  // 32'hf36448a0;
    ram_cell[     260] = 32'h0;  // 32'h1a8593fe;
    ram_cell[     261] = 32'h0;  // 32'h633c8349;
    ram_cell[     262] = 32'h0;  // 32'h508ebe61;
    ram_cell[     263] = 32'h0;  // 32'hef3d108b;
    ram_cell[     264] = 32'h0;  // 32'hc44bdd4e;
    ram_cell[     265] = 32'h0;  // 32'hcccf3dfa;
    ram_cell[     266] = 32'h0;  // 32'h81bcb0aa;
    ram_cell[     267] = 32'h0;  // 32'h7a24cdf3;
    ram_cell[     268] = 32'h0;  // 32'hff664800;
    ram_cell[     269] = 32'h0;  // 32'h04c4332b;
    ram_cell[     270] = 32'h0;  // 32'h339b3764;
    ram_cell[     271] = 32'h0;  // 32'h30f9b303;
    ram_cell[     272] = 32'h0;  // 32'h06e8913e;
    ram_cell[     273] = 32'h0;  // 32'ha65e50aa;
    ram_cell[     274] = 32'h0;  // 32'hbef18197;
    ram_cell[     275] = 32'h0;  // 32'ha0c17ca9;
    ram_cell[     276] = 32'h0;  // 32'hdd8b54ed;
    ram_cell[     277] = 32'h0;  // 32'h2ca90cd8;
    ram_cell[     278] = 32'h0;  // 32'h6c5c26eb;
    ram_cell[     279] = 32'h0;  // 32'h63c138ac;
    ram_cell[     280] = 32'h0;  // 32'hff374529;
    ram_cell[     281] = 32'h0;  // 32'h6eb3045f;
    ram_cell[     282] = 32'h0;  // 32'h54d3df46;
    ram_cell[     283] = 32'h0;  // 32'he118f106;
    ram_cell[     284] = 32'h0;  // 32'hf83716b2;
    ram_cell[     285] = 32'h0;  // 32'hc49a83e9;
    ram_cell[     286] = 32'h0;  // 32'hafc3c730;
    ram_cell[     287] = 32'h0;  // 32'hcdd2cabf;
    ram_cell[     288] = 32'h0;  // 32'h2973fa10;
    ram_cell[     289] = 32'h0;  // 32'h8f044b9d;
    ram_cell[     290] = 32'h0;  // 32'he01e0c5e;
    ram_cell[     291] = 32'h0;  // 32'h4b7ddcc6;
    ram_cell[     292] = 32'h0;  // 32'ha91b98d0;
    ram_cell[     293] = 32'h0;  // 32'h971a7160;
    ram_cell[     294] = 32'h0;  // 32'h0e624fc1;
    ram_cell[     295] = 32'h0;  // 32'hc9afed43;
    ram_cell[     296] = 32'h0;  // 32'haba1266a;
    ram_cell[     297] = 32'h0;  // 32'hcb7637a7;
    ram_cell[     298] = 32'h0;  // 32'h42721742;
    ram_cell[     299] = 32'h0;  // 32'hd4a9b095;
    ram_cell[     300] = 32'h0;  // 32'h0ef3f824;
    ram_cell[     301] = 32'h0;  // 32'h978607a3;
    ram_cell[     302] = 32'h0;  // 32'h8ae85e8e;
    ram_cell[     303] = 32'h0;  // 32'h1c5c9504;
    ram_cell[     304] = 32'h0;  // 32'h90767897;
    ram_cell[     305] = 32'h0;  // 32'h2a773baa;
    ram_cell[     306] = 32'h0;  // 32'h220ae560;
    ram_cell[     307] = 32'h0;  // 32'he27e28fb;
    ram_cell[     308] = 32'h0;  // 32'hbe91ec9a;
    ram_cell[     309] = 32'h0;  // 32'h91483afc;
    ram_cell[     310] = 32'h0;  // 32'h80fe4702;
    ram_cell[     311] = 32'h0;  // 32'h4a0a9185;
    ram_cell[     312] = 32'h0;  // 32'hd2ca7578;
    ram_cell[     313] = 32'h0;  // 32'he27090bd;
    ram_cell[     314] = 32'h0;  // 32'hdb765d64;
    ram_cell[     315] = 32'h0;  // 32'h3d8bfb50;
    ram_cell[     316] = 32'h0;  // 32'hc9bc4c08;
    ram_cell[     317] = 32'h0;  // 32'hb948eff3;
    ram_cell[     318] = 32'h0;  // 32'h64194c2a;
    ram_cell[     319] = 32'h0;  // 32'hb743a8c8;
    ram_cell[     320] = 32'h0;  // 32'h80d9a2e0;
    ram_cell[     321] = 32'h0;  // 32'h42efe98e;
    ram_cell[     322] = 32'h0;  // 32'h7c26234e;
    ram_cell[     323] = 32'h0;  // 32'h8234ee0f;
    ram_cell[     324] = 32'h0;  // 32'h898f92f5;
    ram_cell[     325] = 32'h0;  // 32'h7a9a4edf;
    ram_cell[     326] = 32'h0;  // 32'h350e324a;
    ram_cell[     327] = 32'h0;  // 32'h5130c96a;
    ram_cell[     328] = 32'h0;  // 32'h16c3cb39;
    ram_cell[     329] = 32'h0;  // 32'hf2e8049c;
    ram_cell[     330] = 32'h0;  // 32'h2e3e33ef;
    ram_cell[     331] = 32'h0;  // 32'h6c1fcd61;
    ram_cell[     332] = 32'h0;  // 32'h9a294356;
    ram_cell[     333] = 32'h0;  // 32'hcae4e6d0;
    ram_cell[     334] = 32'h0;  // 32'h9b044c09;
    ram_cell[     335] = 32'h0;  // 32'h1cc28578;
    ram_cell[     336] = 32'h0;  // 32'h2d99fa6c;
    ram_cell[     337] = 32'h0;  // 32'hbcd06308;
    ram_cell[     338] = 32'h0;  // 32'h4888158e;
    ram_cell[     339] = 32'h0;  // 32'h2180c306;
    ram_cell[     340] = 32'h0;  // 32'h633d194c;
    ram_cell[     341] = 32'h0;  // 32'hd44b521b;
    ram_cell[     342] = 32'h0;  // 32'h8e70a08a;
    ram_cell[     343] = 32'h0;  // 32'ha67e3174;
    ram_cell[     344] = 32'h0;  // 32'h59e62bf8;
    ram_cell[     345] = 32'h0;  // 32'h95d89d73;
    ram_cell[     346] = 32'h0;  // 32'hf63c3517;
    ram_cell[     347] = 32'h0;  // 32'hebdf0f66;
    ram_cell[     348] = 32'h0;  // 32'he93c4c8c;
    ram_cell[     349] = 32'h0;  // 32'ha5be53e1;
    ram_cell[     350] = 32'h0;  // 32'h659c806c;
    ram_cell[     351] = 32'h0;  // 32'h0d4afe2f;
    ram_cell[     352] = 32'h0;  // 32'hf1e7f50d;
    ram_cell[     353] = 32'h0;  // 32'hadfce948;
    ram_cell[     354] = 32'h0;  // 32'hc8b552b7;
    ram_cell[     355] = 32'h0;  // 32'hc435b0a8;
    ram_cell[     356] = 32'h0;  // 32'h938956e4;
    ram_cell[     357] = 32'h0;  // 32'h4f90e78a;
    ram_cell[     358] = 32'h0;  // 32'h06665e85;
    ram_cell[     359] = 32'h0;  // 32'h083d73df;
    ram_cell[     360] = 32'h0;  // 32'h62b4bf23;
    ram_cell[     361] = 32'h0;  // 32'hac963d53;
    ram_cell[     362] = 32'h0;  // 32'h95e6b96c;
    ram_cell[     363] = 32'h0;  // 32'h90e59f24;
    ram_cell[     364] = 32'h0;  // 32'hbcfbc7a8;
    ram_cell[     365] = 32'h0;  // 32'hdc94c25d;
    ram_cell[     366] = 32'h0;  // 32'ha0b348be;
    ram_cell[     367] = 32'h0;  // 32'hb0a3f2c5;
    ram_cell[     368] = 32'h0;  // 32'h6618849d;
    ram_cell[     369] = 32'h0;  // 32'h43109a43;
    ram_cell[     370] = 32'h0;  // 32'hbf8e3e55;
    ram_cell[     371] = 32'h0;  // 32'h13a1b140;
    ram_cell[     372] = 32'h0;  // 32'he26a5ca0;
    ram_cell[     373] = 32'h0;  // 32'h8ba43cf9;
    ram_cell[     374] = 32'h0;  // 32'he7a20939;
    ram_cell[     375] = 32'h0;  // 32'h8eb8aea6;
    ram_cell[     376] = 32'h0;  // 32'he526d6b0;
    ram_cell[     377] = 32'h0;  // 32'h6ae81f4b;
    ram_cell[     378] = 32'h0;  // 32'hd828cb1b;
    ram_cell[     379] = 32'h0;  // 32'he9c5388b;
    ram_cell[     380] = 32'h0;  // 32'h158ce910;
    ram_cell[     381] = 32'h0;  // 32'he2bf3586;
    ram_cell[     382] = 32'h0;  // 32'h9150caa0;
    ram_cell[     383] = 32'h0;  // 32'h8cc1cdf1;
    ram_cell[     384] = 32'h0;  // 32'h24b58efb;
    ram_cell[     385] = 32'h0;  // 32'h610412a4;
    ram_cell[     386] = 32'h0;  // 32'he90bf2cd;
    ram_cell[     387] = 32'h0;  // 32'ha23bdc45;
    ram_cell[     388] = 32'h0;  // 32'hec7354ba;
    ram_cell[     389] = 32'h0;  // 32'h61a680a9;
    ram_cell[     390] = 32'h0;  // 32'hee91855c;
    ram_cell[     391] = 32'h0;  // 32'hc8caab1d;
    ram_cell[     392] = 32'h0;  // 32'h6effba14;
    ram_cell[     393] = 32'h0;  // 32'h068ea1e9;
    ram_cell[     394] = 32'h0;  // 32'hb7fca25c;
    ram_cell[     395] = 32'h0;  // 32'h7d81945e;
    ram_cell[     396] = 32'h0;  // 32'h1735f559;
    ram_cell[     397] = 32'h0;  // 32'h5973ff1b;
    ram_cell[     398] = 32'h0;  // 32'h84f943f6;
    ram_cell[     399] = 32'h0;  // 32'h31b4ef31;
    ram_cell[     400] = 32'h0;  // 32'ha064781d;
    ram_cell[     401] = 32'h0;  // 32'he9fc11cb;
    ram_cell[     402] = 32'h0;  // 32'h7145b6d1;
    ram_cell[     403] = 32'h0;  // 32'hc8b98fc3;
    ram_cell[     404] = 32'h0;  // 32'h96838286;
    ram_cell[     405] = 32'h0;  // 32'hb855b928;
    ram_cell[     406] = 32'h0;  // 32'h36db87d6;
    ram_cell[     407] = 32'h0;  // 32'h7428161a;
    ram_cell[     408] = 32'h0;  // 32'hb64f82d3;
    ram_cell[     409] = 32'h0;  // 32'h429137b9;
    ram_cell[     410] = 32'h0;  // 32'h45ab8095;
    ram_cell[     411] = 32'h0;  // 32'h8376d415;
    ram_cell[     412] = 32'h0;  // 32'h9aa72f6b;
    ram_cell[     413] = 32'h0;  // 32'h90db7741;
    ram_cell[     414] = 32'h0;  // 32'h1bf04433;
    ram_cell[     415] = 32'h0;  // 32'hb1c2c9b7;
    ram_cell[     416] = 32'h0;  // 32'h495ab4cf;
    ram_cell[     417] = 32'h0;  // 32'h55ab13cb;
    ram_cell[     418] = 32'h0;  // 32'hbc2afd8a;
    ram_cell[     419] = 32'h0;  // 32'hec1b1344;
    ram_cell[     420] = 32'h0;  // 32'h5c0e49cf;
    ram_cell[     421] = 32'h0;  // 32'hf052aa26;
    ram_cell[     422] = 32'h0;  // 32'haabe8bf8;
    ram_cell[     423] = 32'h0;  // 32'h81ee6427;
    ram_cell[     424] = 32'h0;  // 32'hde5282ae;
    ram_cell[     425] = 32'h0;  // 32'h0aa934bc;
    ram_cell[     426] = 32'h0;  // 32'hb582a735;
    ram_cell[     427] = 32'h0;  // 32'h44e6af4f;
    ram_cell[     428] = 32'h0;  // 32'hc36021f3;
    ram_cell[     429] = 32'h0;  // 32'hdfd95f3b;
    ram_cell[     430] = 32'h0;  // 32'h54b35121;
    ram_cell[     431] = 32'h0;  // 32'h5c4bd9d7;
    ram_cell[     432] = 32'h0;  // 32'h54abfe92;
    ram_cell[     433] = 32'h0;  // 32'h017d5786;
    ram_cell[     434] = 32'h0;  // 32'hb739c30a;
    ram_cell[     435] = 32'h0;  // 32'h6387e864;
    ram_cell[     436] = 32'h0;  // 32'h77653ad0;
    ram_cell[     437] = 32'h0;  // 32'h7506ef40;
    ram_cell[     438] = 32'h0;  // 32'h25583a25;
    ram_cell[     439] = 32'h0;  // 32'h8106b506;
    ram_cell[     440] = 32'h0;  // 32'he9a91423;
    ram_cell[     441] = 32'h0;  // 32'h93de4a12;
    ram_cell[     442] = 32'h0;  // 32'h608a0af6;
    ram_cell[     443] = 32'h0;  // 32'h0d7049fa;
    ram_cell[     444] = 32'h0;  // 32'h8f32bc08;
    ram_cell[     445] = 32'h0;  // 32'h628a46e8;
    ram_cell[     446] = 32'h0;  // 32'h46452bc2;
    ram_cell[     447] = 32'h0;  // 32'h5ee5c604;
    ram_cell[     448] = 32'h0;  // 32'hd16d1479;
    ram_cell[     449] = 32'h0;  // 32'h3c5184d8;
    ram_cell[     450] = 32'h0;  // 32'hb67a9e25;
    ram_cell[     451] = 32'h0;  // 32'h160a828f;
    ram_cell[     452] = 32'h0;  // 32'h25e0823c;
    ram_cell[     453] = 32'h0;  // 32'hc625b004;
    ram_cell[     454] = 32'h0;  // 32'h5b811a2a;
    ram_cell[     455] = 32'h0;  // 32'ha45551b8;
    ram_cell[     456] = 32'h0;  // 32'hd37c7f8a;
    ram_cell[     457] = 32'h0;  // 32'ha61e48fb;
    ram_cell[     458] = 32'h0;  // 32'h2212edf0;
    ram_cell[     459] = 32'h0;  // 32'h2dd46cdf;
    ram_cell[     460] = 32'h0;  // 32'h3d74c55e;
    ram_cell[     461] = 32'h0;  // 32'h3dafffbd;
    ram_cell[     462] = 32'h0;  // 32'hd3ecfa8b;
    ram_cell[     463] = 32'h0;  // 32'ha6f65d51;
    ram_cell[     464] = 32'h0;  // 32'hfe42854d;
    ram_cell[     465] = 32'h0;  // 32'ha2ffdfd3;
    ram_cell[     466] = 32'h0;  // 32'hfff42d84;
    ram_cell[     467] = 32'h0;  // 32'hefb08b7c;
    ram_cell[     468] = 32'h0;  // 32'h1e7a7e61;
    ram_cell[     469] = 32'h0;  // 32'hd5ec9ef5;
    ram_cell[     470] = 32'h0;  // 32'hdd59b54f;
    ram_cell[     471] = 32'h0;  // 32'h0f396772;
    ram_cell[     472] = 32'h0;  // 32'h9c86d055;
    ram_cell[     473] = 32'h0;  // 32'hb48b0a69;
    ram_cell[     474] = 32'h0;  // 32'h959c83b5;
    ram_cell[     475] = 32'h0;  // 32'hbd69a9c5;
    ram_cell[     476] = 32'h0;  // 32'hcf4468d9;
    ram_cell[     477] = 32'h0;  // 32'h3908d8ae;
    ram_cell[     478] = 32'h0;  // 32'h821bada9;
    ram_cell[     479] = 32'h0;  // 32'h5e5005c1;
    ram_cell[     480] = 32'h0;  // 32'habf73c31;
    ram_cell[     481] = 32'h0;  // 32'h424f999b;
    ram_cell[     482] = 32'h0;  // 32'he47e5143;
    ram_cell[     483] = 32'h0;  // 32'h576571af;
    ram_cell[     484] = 32'h0;  // 32'h90875d74;
    ram_cell[     485] = 32'h0;  // 32'h22ce4348;
    ram_cell[     486] = 32'h0;  // 32'h982ff942;
    ram_cell[     487] = 32'h0;  // 32'hb5063461;
    ram_cell[     488] = 32'h0;  // 32'hb855ac25;
    ram_cell[     489] = 32'h0;  // 32'hc621d5b9;
    ram_cell[     490] = 32'h0;  // 32'h0f1f95bb;
    ram_cell[     491] = 32'h0;  // 32'h3e15f926;
    ram_cell[     492] = 32'h0;  // 32'h771d4016;
    ram_cell[     493] = 32'h0;  // 32'hd24775f6;
    ram_cell[     494] = 32'h0;  // 32'h76a43a9f;
    ram_cell[     495] = 32'h0;  // 32'h7af2659e;
    ram_cell[     496] = 32'h0;  // 32'h960f4554;
    ram_cell[     497] = 32'h0;  // 32'h439a0f12;
    ram_cell[     498] = 32'h0;  // 32'hf8eda8de;
    ram_cell[     499] = 32'h0;  // 32'h337085a9;
    ram_cell[     500] = 32'h0;  // 32'h6c7fb59a;
    ram_cell[     501] = 32'h0;  // 32'he2fe5128;
    ram_cell[     502] = 32'h0;  // 32'he03b4aa6;
    ram_cell[     503] = 32'h0;  // 32'h3d21b46e;
    ram_cell[     504] = 32'h0;  // 32'h9b1ace8e;
    ram_cell[     505] = 32'h0;  // 32'h33306c7b;
    ram_cell[     506] = 32'h0;  // 32'h5ba085de;
    ram_cell[     507] = 32'h0;  // 32'h7a0a2cf0;
    ram_cell[     508] = 32'h0;  // 32'h5118b81c;
    ram_cell[     509] = 32'h0;  // 32'hdae715a5;
    ram_cell[     510] = 32'h0;  // 32'h317993ed;
    ram_cell[     511] = 32'h0;  // 32'h9abc60f9;
    ram_cell[     512] = 32'h0;  // 32'h1b4b5b2b;
    ram_cell[     513] = 32'h0;  // 32'he4d0580c;
    ram_cell[     514] = 32'h0;  // 32'h8eef1946;
    ram_cell[     515] = 32'h0;  // 32'hccb7c2f5;
    ram_cell[     516] = 32'h0;  // 32'h456be70e;
    ram_cell[     517] = 32'h0;  // 32'h8eaec21e;
    ram_cell[     518] = 32'h0;  // 32'hfc05428a;
    ram_cell[     519] = 32'h0;  // 32'h38ad096e;
    ram_cell[     520] = 32'h0;  // 32'h8e70407b;
    ram_cell[     521] = 32'h0;  // 32'hbca5019a;
    ram_cell[     522] = 32'h0;  // 32'h8896396a;
    ram_cell[     523] = 32'h0;  // 32'h157e0c44;
    ram_cell[     524] = 32'h0;  // 32'h673cc08f;
    ram_cell[     525] = 32'h0;  // 32'h1d16a8ba;
    ram_cell[     526] = 32'h0;  // 32'h6829f90c;
    ram_cell[     527] = 32'h0;  // 32'h694d6a65;
    ram_cell[     528] = 32'h0;  // 32'hf598636f;
    ram_cell[     529] = 32'h0;  // 32'h8d34523e;
    ram_cell[     530] = 32'h0;  // 32'h1066c764;
    ram_cell[     531] = 32'h0;  // 32'h7b6dbb27;
    ram_cell[     532] = 32'h0;  // 32'h2bfc4bbd;
    ram_cell[     533] = 32'h0;  // 32'h2e4dc0b2;
    ram_cell[     534] = 32'h0;  // 32'he43c830c;
    ram_cell[     535] = 32'h0;  // 32'h81133a53;
    ram_cell[     536] = 32'h0;  // 32'h48d226a6;
    ram_cell[     537] = 32'h0;  // 32'h2c945fb1;
    ram_cell[     538] = 32'h0;  // 32'hdeae7d8d;
    ram_cell[     539] = 32'h0;  // 32'h12b335a0;
    ram_cell[     540] = 32'h0;  // 32'hf5e1dc53;
    ram_cell[     541] = 32'h0;  // 32'hf6eb4b89;
    ram_cell[     542] = 32'h0;  // 32'h5e5a8b58;
    ram_cell[     543] = 32'h0;  // 32'h951558d8;
    ram_cell[     544] = 32'h0;  // 32'he93d6716;
    ram_cell[     545] = 32'h0;  // 32'hb09cad11;
    ram_cell[     546] = 32'h0;  // 32'h9d2f2f67;
    ram_cell[     547] = 32'h0;  // 32'ha67c891a;
    ram_cell[     548] = 32'h0;  // 32'ha941b279;
    ram_cell[     549] = 32'h0;  // 32'h3349f1e5;
    ram_cell[     550] = 32'h0;  // 32'hd5d934e3;
    ram_cell[     551] = 32'h0;  // 32'h6bb2902f;
    ram_cell[     552] = 32'h0;  // 32'hed7a41d3;
    ram_cell[     553] = 32'h0;  // 32'hc550663e;
    ram_cell[     554] = 32'h0;  // 32'h2a7af8ff;
    ram_cell[     555] = 32'h0;  // 32'h1e77ffe9;
    ram_cell[     556] = 32'h0;  // 32'h44afcfe9;
    ram_cell[     557] = 32'h0;  // 32'h6e34c167;
    ram_cell[     558] = 32'h0;  // 32'ha1546a40;
    ram_cell[     559] = 32'h0;  // 32'h6d2e9cf1;
    ram_cell[     560] = 32'h0;  // 32'hf0ce0990;
    ram_cell[     561] = 32'h0;  // 32'h740ff24c;
    ram_cell[     562] = 32'h0;  // 32'hbe1a7a98;
    ram_cell[     563] = 32'h0;  // 32'h717f9feb;
    ram_cell[     564] = 32'h0;  // 32'hf01f965e;
    ram_cell[     565] = 32'h0;  // 32'hb306772e;
    ram_cell[     566] = 32'h0;  // 32'hfe0a2cdb;
    ram_cell[     567] = 32'h0;  // 32'hbb4c1bbb;
    ram_cell[     568] = 32'h0;  // 32'h6fb72d1f;
    ram_cell[     569] = 32'h0;  // 32'h2fd07a1e;
    ram_cell[     570] = 32'h0;  // 32'h44ac2bf4;
    ram_cell[     571] = 32'h0;  // 32'h0b55406c;
    ram_cell[     572] = 32'h0;  // 32'h64e4dabb;
    ram_cell[     573] = 32'h0;  // 32'h77c256c0;
    ram_cell[     574] = 32'h0;  // 32'h9d136b2a;
    ram_cell[     575] = 32'h0;  // 32'h592ba92e;
    ram_cell[     576] = 32'h0;  // 32'hf9f6d528;
    ram_cell[     577] = 32'h0;  // 32'h9c33366b;
    ram_cell[     578] = 32'h0;  // 32'hf517a756;
    ram_cell[     579] = 32'h0;  // 32'h7d213851;
    ram_cell[     580] = 32'h0;  // 32'h901c1f0d;
    ram_cell[     581] = 32'h0;  // 32'h1bceba6f;
    ram_cell[     582] = 32'h0;  // 32'h5e10e289;
    ram_cell[     583] = 32'h0;  // 32'h6b86d8ef;
    ram_cell[     584] = 32'h0;  // 32'hf12769ce;
    ram_cell[     585] = 32'h0;  // 32'ha2e038c7;
    ram_cell[     586] = 32'h0;  // 32'h9567b5aa;
    ram_cell[     587] = 32'h0;  // 32'ha00b98f8;
    ram_cell[     588] = 32'h0;  // 32'h55caf89c;
    ram_cell[     589] = 32'h0;  // 32'he9b97f16;
    ram_cell[     590] = 32'h0;  // 32'h7c4f98a5;
    ram_cell[     591] = 32'h0;  // 32'h537238d8;
    ram_cell[     592] = 32'h0;  // 32'hb381cdbc;
    ram_cell[     593] = 32'h0;  // 32'he0aa244d;
    ram_cell[     594] = 32'h0;  // 32'h5bd080c7;
    ram_cell[     595] = 32'h0;  // 32'h9713fc5b;
    ram_cell[     596] = 32'h0;  // 32'h7f74736f;
    ram_cell[     597] = 32'h0;  // 32'hec19252d;
    ram_cell[     598] = 32'h0;  // 32'h24fca8e4;
    ram_cell[     599] = 32'h0;  // 32'hd5037472;
    ram_cell[     600] = 32'h0;  // 32'h7d3222b8;
    ram_cell[     601] = 32'h0;  // 32'h00b7e063;
    ram_cell[     602] = 32'h0;  // 32'h20b56554;
    ram_cell[     603] = 32'h0;  // 32'h74bb9f53;
    ram_cell[     604] = 32'h0;  // 32'h9ed647e8;
    ram_cell[     605] = 32'h0;  // 32'hd5180dbc;
    ram_cell[     606] = 32'h0;  // 32'h6725af22;
    ram_cell[     607] = 32'h0;  // 32'hadc6950e;
    ram_cell[     608] = 32'h0;  // 32'hfd58dd52;
    ram_cell[     609] = 32'h0;  // 32'hc91ee775;
    ram_cell[     610] = 32'h0;  // 32'h82905f42;
    ram_cell[     611] = 32'h0;  // 32'h599a681d;
    ram_cell[     612] = 32'h0;  // 32'h6f1dd009;
    ram_cell[     613] = 32'h0;  // 32'h920852a9;
    ram_cell[     614] = 32'h0;  // 32'h55fbc677;
    ram_cell[     615] = 32'h0;  // 32'hd32a1a0a;
    ram_cell[     616] = 32'h0;  // 32'h8e1cf8a3;
    ram_cell[     617] = 32'h0;  // 32'h4c654da4;
    ram_cell[     618] = 32'h0;  // 32'he4ffddd1;
    ram_cell[     619] = 32'h0;  // 32'h6326cb6f;
    ram_cell[     620] = 32'h0;  // 32'h52fa17ff;
    ram_cell[     621] = 32'h0;  // 32'he22626cd;
    ram_cell[     622] = 32'h0;  // 32'h6569ca41;
    ram_cell[     623] = 32'h0;  // 32'h7e1ca77d;
    ram_cell[     624] = 32'h0;  // 32'h997bb4f9;
    ram_cell[     625] = 32'h0;  // 32'hcaf8fd16;
    ram_cell[     626] = 32'h0;  // 32'hf4c12752;
    ram_cell[     627] = 32'h0;  // 32'h6c48647d;
    ram_cell[     628] = 32'h0;  // 32'h3baf2e00;
    ram_cell[     629] = 32'h0;  // 32'h20d37836;
    ram_cell[     630] = 32'h0;  // 32'he7b91907;
    ram_cell[     631] = 32'h0;  // 32'hf48a5b44;
    ram_cell[     632] = 32'h0;  // 32'hc46a03dc;
    ram_cell[     633] = 32'h0;  // 32'hee9a5dbf;
    ram_cell[     634] = 32'h0;  // 32'h06690b64;
    ram_cell[     635] = 32'h0;  // 32'hd0b40016;
    ram_cell[     636] = 32'h0;  // 32'h03ca1441;
    ram_cell[     637] = 32'h0;  // 32'h9b767f98;
    ram_cell[     638] = 32'h0;  // 32'ha21868e1;
    ram_cell[     639] = 32'h0;  // 32'hc8238213;
    ram_cell[     640] = 32'h0;  // 32'hf6922a35;
    ram_cell[     641] = 32'h0;  // 32'hd4d9c9a7;
    ram_cell[     642] = 32'h0;  // 32'h2286d322;
    ram_cell[     643] = 32'h0;  // 32'hd5aa3966;
    ram_cell[     644] = 32'h0;  // 32'h8481e87b;
    ram_cell[     645] = 32'h0;  // 32'h7877c7cb;
    ram_cell[     646] = 32'h0;  // 32'h10486cfd;
    ram_cell[     647] = 32'h0;  // 32'h9428926e;
    ram_cell[     648] = 32'h0;  // 32'h34503a47;
    ram_cell[     649] = 32'h0;  // 32'hc1bcbc35;
    ram_cell[     650] = 32'h0;  // 32'hae6db63e;
    ram_cell[     651] = 32'h0;  // 32'h520e4b2a;
    ram_cell[     652] = 32'h0;  // 32'h0d70c37b;
    ram_cell[     653] = 32'h0;  // 32'hcbfe82a0;
    ram_cell[     654] = 32'h0;  // 32'h39a276b1;
    ram_cell[     655] = 32'h0;  // 32'hf43d50df;
    ram_cell[     656] = 32'h0;  // 32'h93fb4798;
    ram_cell[     657] = 32'h0;  // 32'ha25062d1;
    ram_cell[     658] = 32'h0;  // 32'h6e5711f6;
    ram_cell[     659] = 32'h0;  // 32'hd4dae5cf;
    ram_cell[     660] = 32'h0;  // 32'hc069ac7a;
    ram_cell[     661] = 32'h0;  // 32'h307a6575;
    ram_cell[     662] = 32'h0;  // 32'h019288b3;
    ram_cell[     663] = 32'h0;  // 32'h269b3fac;
    ram_cell[     664] = 32'h0;  // 32'he5e710ac;
    ram_cell[     665] = 32'h0;  // 32'h098c2d5a;
    ram_cell[     666] = 32'h0;  // 32'h457add90;
    ram_cell[     667] = 32'h0;  // 32'ha0eccf9b;
    ram_cell[     668] = 32'h0;  // 32'hf67b5890;
    ram_cell[     669] = 32'h0;  // 32'h0b816d32;
    ram_cell[     670] = 32'h0;  // 32'h501193f0;
    ram_cell[     671] = 32'h0;  // 32'he6b1c329;
    ram_cell[     672] = 32'h0;  // 32'hc99d6a07;
    ram_cell[     673] = 32'h0;  // 32'h351d206a;
    ram_cell[     674] = 32'h0;  // 32'hecf8168c;
    ram_cell[     675] = 32'h0;  // 32'h757340e7;
    ram_cell[     676] = 32'h0;  // 32'h058d73e5;
    ram_cell[     677] = 32'h0;  // 32'h0f68ce53;
    ram_cell[     678] = 32'h0;  // 32'he5254240;
    ram_cell[     679] = 32'h0;  // 32'h0bb7e4f4;
    ram_cell[     680] = 32'h0;  // 32'h68380188;
    ram_cell[     681] = 32'h0;  // 32'h35376dd4;
    ram_cell[     682] = 32'h0;  // 32'h35528f6f;
    ram_cell[     683] = 32'h0;  // 32'haa2de585;
    ram_cell[     684] = 32'h0;  // 32'hb3f4cae7;
    ram_cell[     685] = 32'h0;  // 32'ha2dc95de;
    ram_cell[     686] = 32'h0;  // 32'hb9da29bf;
    ram_cell[     687] = 32'h0;  // 32'h058ff216;
    ram_cell[     688] = 32'h0;  // 32'hdad54c37;
    ram_cell[     689] = 32'h0;  // 32'ha6f5c9b1;
    ram_cell[     690] = 32'h0;  // 32'hebc5701b;
    ram_cell[     691] = 32'h0;  // 32'h2932b05e;
    ram_cell[     692] = 32'h0;  // 32'h294e5127;
    ram_cell[     693] = 32'h0;  // 32'h11fd0a8e;
    ram_cell[     694] = 32'h0;  // 32'hc247a411;
    ram_cell[     695] = 32'h0;  // 32'hbb76985b;
    ram_cell[     696] = 32'h0;  // 32'hdbece478;
    ram_cell[     697] = 32'h0;  // 32'h3c5eaaad;
    ram_cell[     698] = 32'h0;  // 32'h926eaeb2;
    ram_cell[     699] = 32'h0;  // 32'h49e89355;
    ram_cell[     700] = 32'h0;  // 32'hae4e9a38;
    ram_cell[     701] = 32'h0;  // 32'h85f359a1;
    ram_cell[     702] = 32'h0;  // 32'hdf791b24;
    ram_cell[     703] = 32'h0;  // 32'hf2468108;
    ram_cell[     704] = 32'h0;  // 32'ha30b180e;
    ram_cell[     705] = 32'h0;  // 32'hbb33ffcc;
    ram_cell[     706] = 32'h0;  // 32'h5f7cf259;
    ram_cell[     707] = 32'h0;  // 32'h60091fc7;
    ram_cell[     708] = 32'h0;  // 32'hf04ef5c3;
    ram_cell[     709] = 32'h0;  // 32'hda7bc1ce;
    ram_cell[     710] = 32'h0;  // 32'hc108d122;
    ram_cell[     711] = 32'h0;  // 32'h3ede69c6;
    ram_cell[     712] = 32'h0;  // 32'h3b5775fa;
    ram_cell[     713] = 32'h0;  // 32'hc3f796b5;
    ram_cell[     714] = 32'h0;  // 32'h8aaa1840;
    ram_cell[     715] = 32'h0;  // 32'h28a0a76f;
    ram_cell[     716] = 32'h0;  // 32'hdafcdea1;
    ram_cell[     717] = 32'h0;  // 32'hcad4ef0b;
    ram_cell[     718] = 32'h0;  // 32'hb24c0ed5;
    ram_cell[     719] = 32'h0;  // 32'h1e7d2f64;
    ram_cell[     720] = 32'h0;  // 32'h528bed17;
    ram_cell[     721] = 32'h0;  // 32'h970051af;
    ram_cell[     722] = 32'h0;  // 32'h7fc0e3f4;
    ram_cell[     723] = 32'h0;  // 32'h00dcc9c6;
    ram_cell[     724] = 32'h0;  // 32'h804d9718;
    ram_cell[     725] = 32'h0;  // 32'h7139375b;
    ram_cell[     726] = 32'h0;  // 32'hb27b8277;
    ram_cell[     727] = 32'h0;  // 32'hd82406f5;
    ram_cell[     728] = 32'h0;  // 32'hb6161174;
    ram_cell[     729] = 32'h0;  // 32'h1b25abbe;
    ram_cell[     730] = 32'h0;  // 32'h7df64d3f;
    ram_cell[     731] = 32'h0;  // 32'h657ff9d2;
    ram_cell[     732] = 32'h0;  // 32'h26027e61;
    ram_cell[     733] = 32'h0;  // 32'h0662a5df;
    ram_cell[     734] = 32'h0;  // 32'h0e4e9fb7;
    ram_cell[     735] = 32'h0;  // 32'h8ac506b9;
    ram_cell[     736] = 32'h0;  // 32'h98df853e;
    ram_cell[     737] = 32'h0;  // 32'h64165c8a;
    ram_cell[     738] = 32'h0;  // 32'h4300d6a8;
    ram_cell[     739] = 32'h0;  // 32'hf6dfe714;
    ram_cell[     740] = 32'h0;  // 32'he1a6af98;
    ram_cell[     741] = 32'h0;  // 32'h377a8a66;
    ram_cell[     742] = 32'h0;  // 32'h9e7c7113;
    ram_cell[     743] = 32'h0;  // 32'he9254444;
    ram_cell[     744] = 32'h0;  // 32'h53caadef;
    ram_cell[     745] = 32'h0;  // 32'hee0401f6;
    ram_cell[     746] = 32'h0;  // 32'h3b6785f8;
    ram_cell[     747] = 32'h0;  // 32'hfcfd8b07;
    ram_cell[     748] = 32'h0;  // 32'h8becef58;
    ram_cell[     749] = 32'h0;  // 32'hed974737;
    ram_cell[     750] = 32'h0;  // 32'hea4eee17;
    ram_cell[     751] = 32'h0;  // 32'h47d0bf32;
    ram_cell[     752] = 32'h0;  // 32'hcdaf0feb;
    ram_cell[     753] = 32'h0;  // 32'h313a689f;
    ram_cell[     754] = 32'h0;  // 32'hebcf0056;
    ram_cell[     755] = 32'h0;  // 32'haead6047;
    ram_cell[     756] = 32'h0;  // 32'hef63028d;
    ram_cell[     757] = 32'h0;  // 32'h670fb2e8;
    ram_cell[     758] = 32'h0;  // 32'h95cce057;
    ram_cell[     759] = 32'h0;  // 32'hf37cf52a;
    ram_cell[     760] = 32'h0;  // 32'h388a6bc5;
    ram_cell[     761] = 32'h0;  // 32'hfad0ad8a;
    ram_cell[     762] = 32'h0;  // 32'h4f10cd10;
    ram_cell[     763] = 32'h0;  // 32'had19454b;
    ram_cell[     764] = 32'h0;  // 32'haac38d01;
    ram_cell[     765] = 32'h0;  // 32'hdce3a632;
    ram_cell[     766] = 32'h0;  // 32'h26ff4e71;
    ram_cell[     767] = 32'h0;  // 32'h903dd392;
    ram_cell[     768] = 32'h0;  // 32'hd40ff3e4;
    ram_cell[     769] = 32'h0;  // 32'hd186a0a0;
    ram_cell[     770] = 32'h0;  // 32'h349a59f3;
    ram_cell[     771] = 32'h0;  // 32'hbeb6bb1f;
    ram_cell[     772] = 32'h0;  // 32'h74568afa;
    ram_cell[     773] = 32'h0;  // 32'h0397fdf6;
    ram_cell[     774] = 32'h0;  // 32'hc28f0943;
    ram_cell[     775] = 32'h0;  // 32'h0795fe4e;
    ram_cell[     776] = 32'h0;  // 32'h9009560b;
    ram_cell[     777] = 32'h0;  // 32'he9dc4ced;
    ram_cell[     778] = 32'h0;  // 32'h08f16d68;
    ram_cell[     779] = 32'h0;  // 32'he2f50b4a;
    ram_cell[     780] = 32'h0;  // 32'hb4c9f2df;
    ram_cell[     781] = 32'h0;  // 32'h4fe21219;
    ram_cell[     782] = 32'h0;  // 32'hf31d7595;
    ram_cell[     783] = 32'h0;  // 32'ha574921d;
    ram_cell[     784] = 32'h0;  // 32'hd7526368;
    ram_cell[     785] = 32'h0;  // 32'h993c9da8;
    ram_cell[     786] = 32'h0;  // 32'h06f9610e;
    ram_cell[     787] = 32'h0;  // 32'h05f387b8;
    ram_cell[     788] = 32'h0;  // 32'h877a10df;
    ram_cell[     789] = 32'h0;  // 32'h4f8e2369;
    ram_cell[     790] = 32'h0;  // 32'h6c47d242;
    ram_cell[     791] = 32'h0;  // 32'h93a1c4f9;
    ram_cell[     792] = 32'h0;  // 32'h738939af;
    ram_cell[     793] = 32'h0;  // 32'h13450f0f;
    ram_cell[     794] = 32'h0;  // 32'h509f9abb;
    ram_cell[     795] = 32'h0;  // 32'h95b276c4;
    ram_cell[     796] = 32'h0;  // 32'h6b34f9b6;
    ram_cell[     797] = 32'h0;  // 32'h2259bc2a;
    ram_cell[     798] = 32'h0;  // 32'h7c9034f4;
    ram_cell[     799] = 32'h0;  // 32'h4eef4420;
    ram_cell[     800] = 32'h0;  // 32'hb8bc2738;
    ram_cell[     801] = 32'h0;  // 32'he6e685e9;
    ram_cell[     802] = 32'h0;  // 32'h4643e71e;
    ram_cell[     803] = 32'h0;  // 32'h1e42b685;
    ram_cell[     804] = 32'h0;  // 32'he2253f70;
    ram_cell[     805] = 32'h0;  // 32'h9d9b68fb;
    ram_cell[     806] = 32'h0;  // 32'hcc98d0f4;
    ram_cell[     807] = 32'h0;  // 32'h0441d38a;
    ram_cell[     808] = 32'h0;  // 32'h4b841cc1;
    ram_cell[     809] = 32'h0;  // 32'ha2ba902e;
    ram_cell[     810] = 32'h0;  // 32'h617d4fc8;
    ram_cell[     811] = 32'h0;  // 32'h7f24fb64;
    ram_cell[     812] = 32'h0;  // 32'hf22b0869;
    ram_cell[     813] = 32'h0;  // 32'hcff7ba5a;
    ram_cell[     814] = 32'h0;  // 32'h822fdbca;
    ram_cell[     815] = 32'h0;  // 32'hbbe2cd5c;
    ram_cell[     816] = 32'h0;  // 32'h73189cd9;
    ram_cell[     817] = 32'h0;  // 32'h126f8fde;
    ram_cell[     818] = 32'h0;  // 32'h6245fe6e;
    ram_cell[     819] = 32'h0;  // 32'hb06354ed;
    ram_cell[     820] = 32'h0;  // 32'h1a6ea48d;
    ram_cell[     821] = 32'h0;  // 32'h969ce4aa;
    ram_cell[     822] = 32'h0;  // 32'hafd2d015;
    ram_cell[     823] = 32'h0;  // 32'ha6eae5ae;
    ram_cell[     824] = 32'h0;  // 32'h32eb5259;
    ram_cell[     825] = 32'h0;  // 32'h75b5e0a4;
    ram_cell[     826] = 32'h0;  // 32'h9230bb4d;
    ram_cell[     827] = 32'h0;  // 32'h19d953ab;
    ram_cell[     828] = 32'h0;  // 32'hcb4cbe10;
    ram_cell[     829] = 32'h0;  // 32'h7cedad87;
    ram_cell[     830] = 32'h0;  // 32'hbaa4a105;
    ram_cell[     831] = 32'h0;  // 32'h1244fccb;
    ram_cell[     832] = 32'h0;  // 32'hf1d486dd;
    ram_cell[     833] = 32'h0;  // 32'he8c3dbae;
    ram_cell[     834] = 32'h0;  // 32'h9345f766;
    ram_cell[     835] = 32'h0;  // 32'h07e01ff5;
    ram_cell[     836] = 32'h0;  // 32'h87cffa2c;
    ram_cell[     837] = 32'h0;  // 32'hc08abfcb;
    ram_cell[     838] = 32'h0;  // 32'hecf42bea;
    ram_cell[     839] = 32'h0;  // 32'h870107b6;
    ram_cell[     840] = 32'h0;  // 32'h2de1c45f;
    ram_cell[     841] = 32'h0;  // 32'h7166fe4f;
    ram_cell[     842] = 32'h0;  // 32'h172cc49a;
    ram_cell[     843] = 32'h0;  // 32'hced4a66d;
    ram_cell[     844] = 32'h0;  // 32'h82b69e05;
    ram_cell[     845] = 32'h0;  // 32'hd06a48d1;
    ram_cell[     846] = 32'h0;  // 32'haad3cecc;
    ram_cell[     847] = 32'h0;  // 32'h866d14b3;
    ram_cell[     848] = 32'h0;  // 32'h6274bd6a;
    ram_cell[     849] = 32'h0;  // 32'h85cbd66f;
    ram_cell[     850] = 32'h0;  // 32'h09764022;
    ram_cell[     851] = 32'h0;  // 32'h7bb20c14;
    ram_cell[     852] = 32'h0;  // 32'hbda40058;
    ram_cell[     853] = 32'h0;  // 32'h1a6927e7;
    ram_cell[     854] = 32'h0;  // 32'h29b3e7ec;
    ram_cell[     855] = 32'h0;  // 32'h2f58aa03;
    ram_cell[     856] = 32'h0;  // 32'hd9f816fb;
    ram_cell[     857] = 32'h0;  // 32'h0188a86e;
    ram_cell[     858] = 32'h0;  // 32'h62607d13;
    ram_cell[     859] = 32'h0;  // 32'hf822c2f0;
    ram_cell[     860] = 32'h0;  // 32'h683620d9;
    ram_cell[     861] = 32'h0;  // 32'h8bca3a89;
    ram_cell[     862] = 32'h0;  // 32'h55b8ff72;
    ram_cell[     863] = 32'h0;  // 32'h54ea915e;
    ram_cell[     864] = 32'h0;  // 32'h67f687a6;
    ram_cell[     865] = 32'h0;  // 32'h3f231983;
    ram_cell[     866] = 32'h0;  // 32'h64ac7635;
    ram_cell[     867] = 32'h0;  // 32'hc6c1796a;
    ram_cell[     868] = 32'h0;  // 32'h83b98cf0;
    ram_cell[     869] = 32'h0;  // 32'hb3dd3013;
    ram_cell[     870] = 32'h0;  // 32'hef65875e;
    ram_cell[     871] = 32'h0;  // 32'h7b3bb034;
    ram_cell[     872] = 32'h0;  // 32'hb1e76b24;
    ram_cell[     873] = 32'h0;  // 32'h77d3d86d;
    ram_cell[     874] = 32'h0;  // 32'hcb99cbab;
    ram_cell[     875] = 32'h0;  // 32'h80a9d5ff;
    ram_cell[     876] = 32'h0;  // 32'h74659914;
    ram_cell[     877] = 32'h0;  // 32'h26bd9493;
    ram_cell[     878] = 32'h0;  // 32'hae845eed;
    ram_cell[     879] = 32'h0;  // 32'hbed36a31;
    ram_cell[     880] = 32'h0;  // 32'h97a176ae;
    ram_cell[     881] = 32'h0;  // 32'h6adafde2;
    ram_cell[     882] = 32'h0;  // 32'h79a7116f;
    ram_cell[     883] = 32'h0;  // 32'habfb91d9;
    ram_cell[     884] = 32'h0;  // 32'hecdb63be;
    ram_cell[     885] = 32'h0;  // 32'h41d562e2;
    ram_cell[     886] = 32'h0;  // 32'hab54f966;
    ram_cell[     887] = 32'h0;  // 32'h33f9662a;
    ram_cell[     888] = 32'h0;  // 32'h841c1795;
    ram_cell[     889] = 32'h0;  // 32'h25716ae7;
    ram_cell[     890] = 32'h0;  // 32'hef49f8a9;
    ram_cell[     891] = 32'h0;  // 32'h90069f2e;
    ram_cell[     892] = 32'h0;  // 32'h0fdea2f1;
    ram_cell[     893] = 32'h0;  // 32'h5df044f9;
    ram_cell[     894] = 32'h0;  // 32'hb057bd69;
    ram_cell[     895] = 32'h0;  // 32'hd0347746;
    ram_cell[     896] = 32'h0;  // 32'h5ab4cef8;
    ram_cell[     897] = 32'h0;  // 32'h096c3c44;
    ram_cell[     898] = 32'h0;  // 32'hba444563;
    ram_cell[     899] = 32'h0;  // 32'h8cce490a;
    ram_cell[     900] = 32'h0;  // 32'h2415b525;
    ram_cell[     901] = 32'h0;  // 32'he4b35a3a;
    ram_cell[     902] = 32'h0;  // 32'ha5dce470;
    ram_cell[     903] = 32'h0;  // 32'ha977b72a;
    ram_cell[     904] = 32'h0;  // 32'hc2a7d8ba;
    ram_cell[     905] = 32'h0;  // 32'h69810c51;
    ram_cell[     906] = 32'h0;  // 32'haaa62b6b;
    ram_cell[     907] = 32'h0;  // 32'h896c13cf;
    ram_cell[     908] = 32'h0;  // 32'h4d2bb2eb;
    ram_cell[     909] = 32'h0;  // 32'had7c0d8c;
    ram_cell[     910] = 32'h0;  // 32'h3f53d675;
    ram_cell[     911] = 32'h0;  // 32'hd91efd56;
    ram_cell[     912] = 32'h0;  // 32'h39f0b20a;
    ram_cell[     913] = 32'h0;  // 32'h44b4b4da;
    ram_cell[     914] = 32'h0;  // 32'h507f9571;
    ram_cell[     915] = 32'h0;  // 32'hdb9c83f5;
    ram_cell[     916] = 32'h0;  // 32'h065cb3f9;
    ram_cell[     917] = 32'h0;  // 32'h439fef37;
    ram_cell[     918] = 32'h0;  // 32'hd2f27177;
    ram_cell[     919] = 32'h0;  // 32'h0a8691de;
    ram_cell[     920] = 32'h0;  // 32'h95c938af;
    ram_cell[     921] = 32'h0;  // 32'h6fdb5d15;
    ram_cell[     922] = 32'h0;  // 32'h3c67d9e8;
    ram_cell[     923] = 32'h0;  // 32'hd52b0c71;
    ram_cell[     924] = 32'h0;  // 32'h1dc5e25c;
    ram_cell[     925] = 32'h0;  // 32'h69e24e7a;
    ram_cell[     926] = 32'h0;  // 32'h200d2b96;
    ram_cell[     927] = 32'h0;  // 32'h451ee24b;
    ram_cell[     928] = 32'h0;  // 32'he53783ac;
    ram_cell[     929] = 32'h0;  // 32'hc12822a5;
    ram_cell[     930] = 32'h0;  // 32'h740bc847;
    ram_cell[     931] = 32'h0;  // 32'h9e779a5f;
    ram_cell[     932] = 32'h0;  // 32'hdfdd180a;
    ram_cell[     933] = 32'h0;  // 32'hca6a519c;
    ram_cell[     934] = 32'h0;  // 32'hc181ad4a;
    ram_cell[     935] = 32'h0;  // 32'hd7406e00;
    ram_cell[     936] = 32'h0;  // 32'h6147feae;
    ram_cell[     937] = 32'h0;  // 32'h3748b710;
    ram_cell[     938] = 32'h0;  // 32'hdd49c0ed;
    ram_cell[     939] = 32'h0;  // 32'h0abd1add;
    ram_cell[     940] = 32'h0;  // 32'hb343550b;
    ram_cell[     941] = 32'h0;  // 32'hc0897b2a;
    ram_cell[     942] = 32'h0;  // 32'h6e425867;
    ram_cell[     943] = 32'h0;  // 32'hbc66e7d7;
    ram_cell[     944] = 32'h0;  // 32'hac1d5198;
    ram_cell[     945] = 32'h0;  // 32'h7502f2b3;
    ram_cell[     946] = 32'h0;  // 32'hce565470;
    ram_cell[     947] = 32'h0;  // 32'h8ae66094;
    ram_cell[     948] = 32'h0;  // 32'h64ae6783;
    ram_cell[     949] = 32'h0;  // 32'h5a865f2c;
    ram_cell[     950] = 32'h0;  // 32'h6a975e8b;
    ram_cell[     951] = 32'h0;  // 32'hc8d9a88a;
    ram_cell[     952] = 32'h0;  // 32'h0833c6a4;
    ram_cell[     953] = 32'h0;  // 32'h9330525e;
    ram_cell[     954] = 32'h0;  // 32'h7100c079;
    ram_cell[     955] = 32'h0;  // 32'hd738d834;
    ram_cell[     956] = 32'h0;  // 32'ha3bee6ba;
    ram_cell[     957] = 32'h0;  // 32'hf042ef47;
    ram_cell[     958] = 32'h0;  // 32'hb7eb3431;
    ram_cell[     959] = 32'h0;  // 32'h484b02f4;
    ram_cell[     960] = 32'h0;  // 32'hdeee54e1;
    ram_cell[     961] = 32'h0;  // 32'hd301b9b9;
    ram_cell[     962] = 32'h0;  // 32'hec084349;
    ram_cell[     963] = 32'h0;  // 32'hff46bbe9;
    ram_cell[     964] = 32'h0;  // 32'h5b5da98a;
    ram_cell[     965] = 32'h0;  // 32'ha3a841da;
    ram_cell[     966] = 32'h0;  // 32'h8e1abe0d;
    ram_cell[     967] = 32'h0;  // 32'h24e8e70e;
    ram_cell[     968] = 32'h0;  // 32'h868bc0f1;
    ram_cell[     969] = 32'h0;  // 32'hb0ae3e08;
    ram_cell[     970] = 32'h0;  // 32'hc58feb2d;
    ram_cell[     971] = 32'h0;  // 32'hdb0728e7;
    ram_cell[     972] = 32'h0;  // 32'h888617f6;
    ram_cell[     973] = 32'h0;  // 32'ha7b07a78;
    ram_cell[     974] = 32'h0;  // 32'h4b6625d4;
    ram_cell[     975] = 32'h0;  // 32'h833ac8e0;
    ram_cell[     976] = 32'h0;  // 32'h93bf02e8;
    ram_cell[     977] = 32'h0;  // 32'h2bb245a7;
    ram_cell[     978] = 32'h0;  // 32'h1fac2802;
    ram_cell[     979] = 32'h0;  // 32'h65da5c43;
    ram_cell[     980] = 32'h0;  // 32'h5553c95e;
    ram_cell[     981] = 32'h0;  // 32'h60099619;
    ram_cell[     982] = 32'h0;  // 32'hf1424cfa;
    ram_cell[     983] = 32'h0;  // 32'h5470077b;
    ram_cell[     984] = 32'h0;  // 32'hbbf406f0;
    ram_cell[     985] = 32'h0;  // 32'he5641961;
    ram_cell[     986] = 32'h0;  // 32'h72505746;
    ram_cell[     987] = 32'h0;  // 32'h048f0b4c;
    ram_cell[     988] = 32'h0;  // 32'h7c68454e;
    ram_cell[     989] = 32'h0;  // 32'h3e90fc44;
    ram_cell[     990] = 32'h0;  // 32'h3a1faa39;
    ram_cell[     991] = 32'h0;  // 32'h85c8d48f;
    ram_cell[     992] = 32'h0;  // 32'hb93f9397;
    ram_cell[     993] = 32'h0;  // 32'h074232dc;
    ram_cell[     994] = 32'h0;  // 32'h6f232b15;
    ram_cell[     995] = 32'h0;  // 32'h5b62e5aa;
    ram_cell[     996] = 32'h0;  // 32'h7b259fec;
    ram_cell[     997] = 32'h0;  // 32'h01407660;
    ram_cell[     998] = 32'h0;  // 32'h44d32fad;
    ram_cell[     999] = 32'h0;  // 32'h01e6ee76;
    ram_cell[    1000] = 32'h0;  // 32'hdd2d1903;
    ram_cell[    1001] = 32'h0;  // 32'h3799451f;
    ram_cell[    1002] = 32'h0;  // 32'h1a85c5e0;
    ram_cell[    1003] = 32'h0;  // 32'h1ebe763d;
    ram_cell[    1004] = 32'h0;  // 32'hdfebeec4;
    ram_cell[    1005] = 32'h0;  // 32'hab0de72b;
    ram_cell[    1006] = 32'h0;  // 32'hbc008797;
    ram_cell[    1007] = 32'h0;  // 32'h0d4a4ece;
    ram_cell[    1008] = 32'h0;  // 32'hb6f69d76;
    ram_cell[    1009] = 32'h0;  // 32'h315a4d9d;
    ram_cell[    1010] = 32'h0;  // 32'he95d71c5;
    ram_cell[    1011] = 32'h0;  // 32'h08c48d9a;
    ram_cell[    1012] = 32'h0;  // 32'ha39f1823;
    ram_cell[    1013] = 32'h0;  // 32'h0a1b0be5;
    ram_cell[    1014] = 32'h0;  // 32'h26d294fd;
    ram_cell[    1015] = 32'h0;  // 32'h9dd1a97a;
    ram_cell[    1016] = 32'h0;  // 32'h7e915eec;
    ram_cell[    1017] = 32'h0;  // 32'h87c963fd;
    ram_cell[    1018] = 32'h0;  // 32'h78801882;
    ram_cell[    1019] = 32'h0;  // 32'h1c855c71;
    ram_cell[    1020] = 32'h0;  // 32'h01989261;
    ram_cell[    1021] = 32'h0;  // 32'had794836;
    ram_cell[    1022] = 32'h0;  // 32'h8e5a3dad;
    ram_cell[    1023] = 32'h0;  // 32'hc30d4530;
    ram_cell[    1024] = 32'h0;  // 32'hb72d14bd;
    ram_cell[    1025] = 32'h0;  // 32'h712d9ad5;
    ram_cell[    1026] = 32'h0;  // 32'h0a75410b;
    ram_cell[    1027] = 32'h0;  // 32'h0fc35da7;
    ram_cell[    1028] = 32'h0;  // 32'he747f782;
    ram_cell[    1029] = 32'h0;  // 32'h62afd551;
    ram_cell[    1030] = 32'h0;  // 32'hd034f66f;
    ram_cell[    1031] = 32'h0;  // 32'hacbb1b15;
    ram_cell[    1032] = 32'h0;  // 32'h6f12a9d0;
    ram_cell[    1033] = 32'h0;  // 32'h67b8728d;
    ram_cell[    1034] = 32'h0;  // 32'ha3d1a48a;
    ram_cell[    1035] = 32'h0;  // 32'h05f347cc;
    ram_cell[    1036] = 32'h0;  // 32'h4cac9c2b;
    ram_cell[    1037] = 32'h0;  // 32'h9ccf3d5a;
    ram_cell[    1038] = 32'h0;  // 32'h031e2ef2;
    ram_cell[    1039] = 32'h0;  // 32'h48d4ddd6;
    ram_cell[    1040] = 32'h0;  // 32'h1433028e;
    ram_cell[    1041] = 32'h0;  // 32'h65522978;
    ram_cell[    1042] = 32'h0;  // 32'h987357a0;
    ram_cell[    1043] = 32'h0;  // 32'h96abbd61;
    ram_cell[    1044] = 32'h0;  // 32'hb7a776dd;
    ram_cell[    1045] = 32'h0;  // 32'he860274d;
    ram_cell[    1046] = 32'h0;  // 32'hf94dca44;
    ram_cell[    1047] = 32'h0;  // 32'hc885e580;
    ram_cell[    1048] = 32'h0;  // 32'h2960b85c;
    ram_cell[    1049] = 32'h0;  // 32'h8955edd0;
    ram_cell[    1050] = 32'h0;  // 32'h4325e39e;
    ram_cell[    1051] = 32'h0;  // 32'h1bf5f821;
    ram_cell[    1052] = 32'h0;  // 32'hc453ce45;
    ram_cell[    1053] = 32'h0;  // 32'h0d4682ef;
    ram_cell[    1054] = 32'h0;  // 32'h6723ea47;
    ram_cell[    1055] = 32'h0;  // 32'h6bbb535b;
    ram_cell[    1056] = 32'h0;  // 32'h0cf33f59;
    ram_cell[    1057] = 32'h0;  // 32'ha6526ac7;
    ram_cell[    1058] = 32'h0;  // 32'h9d74ae5e;
    ram_cell[    1059] = 32'h0;  // 32'h119e7d93;
    ram_cell[    1060] = 32'h0;  // 32'h9f8075b9;
    ram_cell[    1061] = 32'h0;  // 32'h1d2436d4;
    ram_cell[    1062] = 32'h0;  // 32'h6dda421e;
    ram_cell[    1063] = 32'h0;  // 32'h3c58d6c8;
    ram_cell[    1064] = 32'h0;  // 32'h7a14c928;
    ram_cell[    1065] = 32'h0;  // 32'h2e4cb7e8;
    ram_cell[    1066] = 32'h0;  // 32'h14081597;
    ram_cell[    1067] = 32'h0;  // 32'hb45668a3;
    ram_cell[    1068] = 32'h0;  // 32'h6847ef1a;
    ram_cell[    1069] = 32'h0;  // 32'hc3c22ab2;
    ram_cell[    1070] = 32'h0;  // 32'h34d98d63;
    ram_cell[    1071] = 32'h0;  // 32'h6fc9f4f8;
    ram_cell[    1072] = 32'h0;  // 32'hbb116b6b;
    ram_cell[    1073] = 32'h0;  // 32'hb4bf9773;
    ram_cell[    1074] = 32'h0;  // 32'h413e4ab0;
    ram_cell[    1075] = 32'h0;  // 32'hb055d7f6;
    ram_cell[    1076] = 32'h0;  // 32'h6f84fa60;
    ram_cell[    1077] = 32'h0;  // 32'h8c8159a0;
    ram_cell[    1078] = 32'h0;  // 32'haceafac1;
    ram_cell[    1079] = 32'h0;  // 32'hf6377a5a;
    ram_cell[    1080] = 32'h0;  // 32'h39a2d18a;
    ram_cell[    1081] = 32'h0;  // 32'h760401de;
    ram_cell[    1082] = 32'h0;  // 32'h76f6a028;
    ram_cell[    1083] = 32'h0;  // 32'h44864c80;
    ram_cell[    1084] = 32'h0;  // 32'hca49ca9d;
    ram_cell[    1085] = 32'h0;  // 32'h2da12413;
    ram_cell[    1086] = 32'h0;  // 32'h87e7aed1;
    ram_cell[    1087] = 32'h0;  // 32'ha5494f13;
    ram_cell[    1088] = 32'h0;  // 32'h7a1fdb4d;
    ram_cell[    1089] = 32'h0;  // 32'h2e310a70;
    ram_cell[    1090] = 32'h0;  // 32'hdb148968;
    ram_cell[    1091] = 32'h0;  // 32'h04afff40;
    ram_cell[    1092] = 32'h0;  // 32'hbfd9316c;
    ram_cell[    1093] = 32'h0;  // 32'h9232c65a;
    ram_cell[    1094] = 32'h0;  // 32'h6d2d5ff1;
    ram_cell[    1095] = 32'h0;  // 32'h7c0b679b;
    ram_cell[    1096] = 32'h0;  // 32'he8502bcc;
    ram_cell[    1097] = 32'h0;  // 32'he3ba1dc2;
    ram_cell[    1098] = 32'h0;  // 32'h5adf57e2;
    ram_cell[    1099] = 32'h0;  // 32'h06a79f56;
    ram_cell[    1100] = 32'h0;  // 32'h14c9f5db;
    ram_cell[    1101] = 32'h0;  // 32'h524381f2;
    ram_cell[    1102] = 32'h0;  // 32'h2c5af4ae;
    ram_cell[    1103] = 32'h0;  // 32'hea0d9023;
    ram_cell[    1104] = 32'h0;  // 32'h95dac484;
    ram_cell[    1105] = 32'h0;  // 32'h77940a5f;
    ram_cell[    1106] = 32'h0;  // 32'h249a7961;
    ram_cell[    1107] = 32'h0;  // 32'h4b87bbd1;
    ram_cell[    1108] = 32'h0;  // 32'h07cda563;
    ram_cell[    1109] = 32'h0;  // 32'h1c30006c;
    ram_cell[    1110] = 32'h0;  // 32'h86fc5227;
    ram_cell[    1111] = 32'h0;  // 32'h5e7e4594;
    ram_cell[    1112] = 32'h0;  // 32'hd7662d72;
    ram_cell[    1113] = 32'h0;  // 32'h67eae660;
    ram_cell[    1114] = 32'h0;  // 32'he0c4ff81;
    ram_cell[    1115] = 32'h0;  // 32'h33ed7f27;
    ram_cell[    1116] = 32'h0;  // 32'hf629683d;
    ram_cell[    1117] = 32'h0;  // 32'hb15bc57b;
    ram_cell[    1118] = 32'h0;  // 32'h1bc3601f;
    ram_cell[    1119] = 32'h0;  // 32'h4f5d7b32;
    ram_cell[    1120] = 32'h0;  // 32'h72869618;
    ram_cell[    1121] = 32'h0;  // 32'hbd890e46;
    ram_cell[    1122] = 32'h0;  // 32'h62039b6f;
    ram_cell[    1123] = 32'h0;  // 32'h88bf1114;
    ram_cell[    1124] = 32'h0;  // 32'ha9332e4f;
    ram_cell[    1125] = 32'h0;  // 32'h97e3b955;
    ram_cell[    1126] = 32'h0;  // 32'h0e0a1bee;
    ram_cell[    1127] = 32'h0;  // 32'h4589126f;
    ram_cell[    1128] = 32'h0;  // 32'hde3c2825;
    ram_cell[    1129] = 32'h0;  // 32'hde074e9f;
    ram_cell[    1130] = 32'h0;  // 32'h5dc5f299;
    ram_cell[    1131] = 32'h0;  // 32'h708f2cd1;
    ram_cell[    1132] = 32'h0;  // 32'h9ecfe83f;
    ram_cell[    1133] = 32'h0;  // 32'hc4aafb3d;
    ram_cell[    1134] = 32'h0;  // 32'ha3d9943e;
    ram_cell[    1135] = 32'h0;  // 32'hd5fb673a;
    ram_cell[    1136] = 32'h0;  // 32'haa9b25af;
    ram_cell[    1137] = 32'h0;  // 32'h8fe9c70f;
    ram_cell[    1138] = 32'h0;  // 32'h3959cc6e;
    ram_cell[    1139] = 32'h0;  // 32'h6c215190;
    ram_cell[    1140] = 32'h0;  // 32'h04cf8b84;
    ram_cell[    1141] = 32'h0;  // 32'hb40de1fb;
    ram_cell[    1142] = 32'h0;  // 32'h370715f2;
    ram_cell[    1143] = 32'h0;  // 32'h0b889c73;
    ram_cell[    1144] = 32'h0;  // 32'hee7d77e3;
    ram_cell[    1145] = 32'h0;  // 32'h333ff63c;
    ram_cell[    1146] = 32'h0;  // 32'h7a8c5019;
    ram_cell[    1147] = 32'h0;  // 32'haa45e8bb;
    ram_cell[    1148] = 32'h0;  // 32'hc38f2401;
    ram_cell[    1149] = 32'h0;  // 32'h38639278;
    ram_cell[    1150] = 32'h0;  // 32'hc8334423;
    ram_cell[    1151] = 32'h0;  // 32'h253a1fdf;
    ram_cell[    1152] = 32'h0;  // 32'h70b4847c;
    ram_cell[    1153] = 32'h0;  // 32'h2c0b7aba;
    ram_cell[    1154] = 32'h0;  // 32'h50ff3a3e;
    ram_cell[    1155] = 32'h0;  // 32'h84c1301d;
    ram_cell[    1156] = 32'h0;  // 32'hcfa9b33e;
    ram_cell[    1157] = 32'h0;  // 32'haa9a73bc;
    ram_cell[    1158] = 32'h0;  // 32'h32ea3a34;
    ram_cell[    1159] = 32'h0;  // 32'haaccb1fe;
    ram_cell[    1160] = 32'h0;  // 32'h5e82b271;
    ram_cell[    1161] = 32'h0;  // 32'h05fb0293;
    ram_cell[    1162] = 32'h0;  // 32'hf924d8bd;
    ram_cell[    1163] = 32'h0;  // 32'hf9a9590a;
    ram_cell[    1164] = 32'h0;  // 32'h06c00135;
    ram_cell[    1165] = 32'h0;  // 32'h4bf8d0db;
    ram_cell[    1166] = 32'h0;  // 32'h2faf198a;
    ram_cell[    1167] = 32'h0;  // 32'h36566aa0;
    ram_cell[    1168] = 32'h0;  // 32'hd27f3fed;
    ram_cell[    1169] = 32'h0;  // 32'hefe0d6fc;
    ram_cell[    1170] = 32'h0;  // 32'hf8dbd6e3;
    ram_cell[    1171] = 32'h0;  // 32'h035accc4;
    ram_cell[    1172] = 32'h0;  // 32'haa3f8e7b;
    ram_cell[    1173] = 32'h0;  // 32'h3bab43c4;
    ram_cell[    1174] = 32'h0;  // 32'h90d10d5e;
    ram_cell[    1175] = 32'h0;  // 32'h05ed5d34;
    ram_cell[    1176] = 32'h0;  // 32'hc8275f75;
    ram_cell[    1177] = 32'h0;  // 32'h0166d884;
    ram_cell[    1178] = 32'h0;  // 32'h9e210e2c;
    ram_cell[    1179] = 32'h0;  // 32'hd3b41ba6;
    ram_cell[    1180] = 32'h0;  // 32'hab67a836;
    ram_cell[    1181] = 32'h0;  // 32'h0914e6cb;
    ram_cell[    1182] = 32'h0;  // 32'h5d904159;
    ram_cell[    1183] = 32'h0;  // 32'hd2fbe820;
    ram_cell[    1184] = 32'h0;  // 32'h5d75d8af;
    ram_cell[    1185] = 32'h0;  // 32'hee516f43;
    ram_cell[    1186] = 32'h0;  // 32'hac07e8ee;
    ram_cell[    1187] = 32'h0;  // 32'h673819e2;
    ram_cell[    1188] = 32'h0;  // 32'h374e9ef4;
    ram_cell[    1189] = 32'h0;  // 32'h5909a4ff;
    ram_cell[    1190] = 32'h0;  // 32'hc4c86e28;
    ram_cell[    1191] = 32'h0;  // 32'hd8dc563b;
    ram_cell[    1192] = 32'h0;  // 32'h512627b8;
    ram_cell[    1193] = 32'h0;  // 32'h650dba93;
    ram_cell[    1194] = 32'h0;  // 32'hdb5c926a;
    ram_cell[    1195] = 32'h0;  // 32'hfbb46000;
    ram_cell[    1196] = 32'h0;  // 32'h0063f7c0;
    ram_cell[    1197] = 32'h0;  // 32'h1690ac4a;
    ram_cell[    1198] = 32'h0;  // 32'h9382fa3f;
    ram_cell[    1199] = 32'h0;  // 32'h98f08cf0;
    ram_cell[    1200] = 32'h0;  // 32'h59a44d37;
    ram_cell[    1201] = 32'h0;  // 32'h24a9f988;
    ram_cell[    1202] = 32'h0;  // 32'h5343f5e8;
    ram_cell[    1203] = 32'h0;  // 32'h019eb8e4;
    ram_cell[    1204] = 32'h0;  // 32'h9c31e4f7;
    ram_cell[    1205] = 32'h0;  // 32'h2f36a403;
    ram_cell[    1206] = 32'h0;  // 32'h6ee8608e;
    ram_cell[    1207] = 32'h0;  // 32'h8dae2a1c;
    ram_cell[    1208] = 32'h0;  // 32'h9092c87b;
    ram_cell[    1209] = 32'h0;  // 32'h88f1818e;
    ram_cell[    1210] = 32'h0;  // 32'hf23b7fe2;
    ram_cell[    1211] = 32'h0;  // 32'hcac651a7;
    ram_cell[    1212] = 32'h0;  // 32'hfaa8c738;
    ram_cell[    1213] = 32'h0;  // 32'hdebf14a7;
    ram_cell[    1214] = 32'h0;  // 32'h620f5628;
    ram_cell[    1215] = 32'h0;  // 32'hee8523fc;
    ram_cell[    1216] = 32'h0;  // 32'hb402d210;
    ram_cell[    1217] = 32'h0;  // 32'he2d55686;
    ram_cell[    1218] = 32'h0;  // 32'h0fcb3978;
    ram_cell[    1219] = 32'h0;  // 32'h75233d88;
    ram_cell[    1220] = 32'h0;  // 32'h0d02495e;
    ram_cell[    1221] = 32'h0;  // 32'h89fe3950;
    ram_cell[    1222] = 32'h0;  // 32'ha34e2158;
    ram_cell[    1223] = 32'h0;  // 32'hb7702916;
    ram_cell[    1224] = 32'h0;  // 32'h30d9b049;
    ram_cell[    1225] = 32'h0;  // 32'h6e0fe32b;
    ram_cell[    1226] = 32'h0;  // 32'h5ef9409a;
    ram_cell[    1227] = 32'h0;  // 32'h39b642a9;
    ram_cell[    1228] = 32'h0;  // 32'hcb2e6aeb;
    ram_cell[    1229] = 32'h0;  // 32'hb5516cc2;
    ram_cell[    1230] = 32'h0;  // 32'h0fdd18fa;
    ram_cell[    1231] = 32'h0;  // 32'hd65e1b23;
    ram_cell[    1232] = 32'h0;  // 32'heeea1116;
    ram_cell[    1233] = 32'h0;  // 32'h81748e35;
    ram_cell[    1234] = 32'h0;  // 32'h6ff0a4cc;
    ram_cell[    1235] = 32'h0;  // 32'h8294873f;
    ram_cell[    1236] = 32'h0;  // 32'h1cab3a24;
    ram_cell[    1237] = 32'h0;  // 32'h394ddb2c;
    ram_cell[    1238] = 32'h0;  // 32'hcc3cdb22;
    ram_cell[    1239] = 32'h0;  // 32'hbd67a79e;
    ram_cell[    1240] = 32'h0;  // 32'h256aa31a;
    ram_cell[    1241] = 32'h0;  // 32'h77df33df;
    ram_cell[    1242] = 32'h0;  // 32'h66052dc1;
    ram_cell[    1243] = 32'h0;  // 32'hfbc08b4d;
    ram_cell[    1244] = 32'h0;  // 32'h56123538;
    ram_cell[    1245] = 32'h0;  // 32'h55833264;
    ram_cell[    1246] = 32'h0;  // 32'h4e0612c0;
    ram_cell[    1247] = 32'h0;  // 32'hd07375e0;
    ram_cell[    1248] = 32'h0;  // 32'hb863acb0;
    ram_cell[    1249] = 32'h0;  // 32'h572f01d3;
    ram_cell[    1250] = 32'h0;  // 32'hf33a6d46;
    ram_cell[    1251] = 32'h0;  // 32'hecd21eb1;
    ram_cell[    1252] = 32'h0;  // 32'h5dbf8e25;
    ram_cell[    1253] = 32'h0;  // 32'h7d32b5ff;
    ram_cell[    1254] = 32'h0;  // 32'h06b9e5f9;
    ram_cell[    1255] = 32'h0;  // 32'h12a81d64;
    ram_cell[    1256] = 32'h0;  // 32'h01b04a30;
    ram_cell[    1257] = 32'h0;  // 32'ha22dcb64;
    ram_cell[    1258] = 32'h0;  // 32'h0278603a;
    ram_cell[    1259] = 32'h0;  // 32'h8d1c3640;
    ram_cell[    1260] = 32'h0;  // 32'h0dad75e1;
    ram_cell[    1261] = 32'h0;  // 32'h0e9282d3;
    ram_cell[    1262] = 32'h0;  // 32'ha6f46a0f;
    ram_cell[    1263] = 32'h0;  // 32'h8485b06b;
    ram_cell[    1264] = 32'h0;  // 32'h15e2cd2c;
    ram_cell[    1265] = 32'h0;  // 32'hfa4b7f45;
    ram_cell[    1266] = 32'h0;  // 32'hbaaf5566;
    ram_cell[    1267] = 32'h0;  // 32'he1ba4cbb;
    ram_cell[    1268] = 32'h0;  // 32'h9a8cda41;
    ram_cell[    1269] = 32'h0;  // 32'habb4dae7;
    ram_cell[    1270] = 32'h0;  // 32'h85f57544;
    ram_cell[    1271] = 32'h0;  // 32'h2cf7d880;
    ram_cell[    1272] = 32'h0;  // 32'h628f1264;
    ram_cell[    1273] = 32'h0;  // 32'hfe2fb072;
    ram_cell[    1274] = 32'h0;  // 32'hc8453f29;
    ram_cell[    1275] = 32'h0;  // 32'h7c6f5950;
    ram_cell[    1276] = 32'h0;  // 32'h70d98cb9;
    ram_cell[    1277] = 32'h0;  // 32'hc163eb3d;
    ram_cell[    1278] = 32'h0;  // 32'h494aae16;
    ram_cell[    1279] = 32'h0;  // 32'h85ccf4c6;
    ram_cell[    1280] = 32'h0;  // 32'hd6a7d1f9;
    ram_cell[    1281] = 32'h0;  // 32'h72f3443e;
    ram_cell[    1282] = 32'h0;  // 32'h8984e615;
    ram_cell[    1283] = 32'h0;  // 32'h4655f3c7;
    ram_cell[    1284] = 32'h0;  // 32'hd8239457;
    ram_cell[    1285] = 32'h0;  // 32'h607d8f29;
    ram_cell[    1286] = 32'h0;  // 32'hb8b85362;
    ram_cell[    1287] = 32'h0;  // 32'h46d67cf3;
    ram_cell[    1288] = 32'h0;  // 32'h7faed202;
    ram_cell[    1289] = 32'h0;  // 32'h695b6f95;
    ram_cell[    1290] = 32'h0;  // 32'h75f11618;
    ram_cell[    1291] = 32'h0;  // 32'h5d72837e;
    ram_cell[    1292] = 32'h0;  // 32'h85924dc2;
    ram_cell[    1293] = 32'h0;  // 32'h31742bef;
    ram_cell[    1294] = 32'h0;  // 32'h6f6c9e01;
    ram_cell[    1295] = 32'h0;  // 32'h6366b05a;
    ram_cell[    1296] = 32'h0;  // 32'h3a321ef2;
    ram_cell[    1297] = 32'h0;  // 32'h202cede3;
    ram_cell[    1298] = 32'h0;  // 32'h907bbc41;
    ram_cell[    1299] = 32'h0;  // 32'h9ecb0272;
    ram_cell[    1300] = 32'h0;  // 32'h63bfc6bd;
    ram_cell[    1301] = 32'h0;  // 32'h27bc1023;
    ram_cell[    1302] = 32'h0;  // 32'h4d2964ca;
    ram_cell[    1303] = 32'h0;  // 32'h57012852;
    ram_cell[    1304] = 32'h0;  // 32'hbe024fa2;
    ram_cell[    1305] = 32'h0;  // 32'h800f7ab8;
    ram_cell[    1306] = 32'h0;  // 32'h1ccdb899;
    ram_cell[    1307] = 32'h0;  // 32'h5daaf1ab;
    ram_cell[    1308] = 32'h0;  // 32'hba690a07;
    ram_cell[    1309] = 32'h0;  // 32'h7b9c79d6;
    ram_cell[    1310] = 32'h0;  // 32'h77e5eb16;
    ram_cell[    1311] = 32'h0;  // 32'h024cf173;
    ram_cell[    1312] = 32'h0;  // 32'hab09a032;
    ram_cell[    1313] = 32'h0;  // 32'h4b93dc45;
    ram_cell[    1314] = 32'h0;  // 32'had5291e9;
    ram_cell[    1315] = 32'h0;  // 32'h65a46fb9;
    ram_cell[    1316] = 32'h0;  // 32'h3e8287c3;
    ram_cell[    1317] = 32'h0;  // 32'hf7312d06;
    ram_cell[    1318] = 32'h0;  // 32'h425c9ded;
    ram_cell[    1319] = 32'h0;  // 32'h82582257;
    ram_cell[    1320] = 32'h0;  // 32'h3f1b0ef7;
    ram_cell[    1321] = 32'h0;  // 32'hb3e9b50a;
    ram_cell[    1322] = 32'h0;  // 32'hbe2e035b;
    ram_cell[    1323] = 32'h0;  // 32'ha5570b95;
    ram_cell[    1324] = 32'h0;  // 32'h2e1f905d;
    ram_cell[    1325] = 32'h0;  // 32'h648a2c4c;
    ram_cell[    1326] = 32'h0;  // 32'h5c961b4a;
    ram_cell[    1327] = 32'h0;  // 32'ha48e6e0f;
    ram_cell[    1328] = 32'h0;  // 32'h52979a0d;
    ram_cell[    1329] = 32'h0;  // 32'h5e19f28f;
    ram_cell[    1330] = 32'h0;  // 32'h29179bbf;
    ram_cell[    1331] = 32'h0;  // 32'h663d7189;
    ram_cell[    1332] = 32'h0;  // 32'h2a34b74d;
    ram_cell[    1333] = 32'h0;  // 32'h943eb458;
    ram_cell[    1334] = 32'h0;  // 32'hb3028fb3;
    ram_cell[    1335] = 32'h0;  // 32'hfbfb71d8;
    ram_cell[    1336] = 32'h0;  // 32'ha725faa9;
    ram_cell[    1337] = 32'h0;  // 32'he035dac2;
    ram_cell[    1338] = 32'h0;  // 32'h615aace3;
    ram_cell[    1339] = 32'h0;  // 32'h5ef0af05;
    ram_cell[    1340] = 32'h0;  // 32'hb425eb0d;
    ram_cell[    1341] = 32'h0;  // 32'hd1fb7e83;
    ram_cell[    1342] = 32'h0;  // 32'hc8f047f9;
    ram_cell[    1343] = 32'h0;  // 32'h41fdfc71;
    ram_cell[    1344] = 32'h0;  // 32'h0a7df7b6;
    ram_cell[    1345] = 32'h0;  // 32'h3469aec6;
    ram_cell[    1346] = 32'h0;  // 32'ha7e0eec3;
    ram_cell[    1347] = 32'h0;  // 32'h11b4f5db;
    ram_cell[    1348] = 32'h0;  // 32'h2c84f81c;
    ram_cell[    1349] = 32'h0;  // 32'h24f88976;
    ram_cell[    1350] = 32'h0;  // 32'h7254df5b;
    ram_cell[    1351] = 32'h0;  // 32'h00021339;
    ram_cell[    1352] = 32'h0;  // 32'h35d30385;
    ram_cell[    1353] = 32'h0;  // 32'h9f94ab94;
    ram_cell[    1354] = 32'h0;  // 32'h604461c9;
    ram_cell[    1355] = 32'h0;  // 32'h90b158a0;
    ram_cell[    1356] = 32'h0;  // 32'h4b06b8fb;
    ram_cell[    1357] = 32'h0;  // 32'hfa26804e;
    ram_cell[    1358] = 32'h0;  // 32'h416c4978;
    ram_cell[    1359] = 32'h0;  // 32'h2589ec42;
    ram_cell[    1360] = 32'h0;  // 32'h20c2a656;
    ram_cell[    1361] = 32'h0;  // 32'h03fab8ce;
    ram_cell[    1362] = 32'h0;  // 32'ha9e17408;
    ram_cell[    1363] = 32'h0;  // 32'h12af5106;
    ram_cell[    1364] = 32'h0;  // 32'h2da57213;
    ram_cell[    1365] = 32'h0;  // 32'hf6fa3341;
    ram_cell[    1366] = 32'h0;  // 32'h75c311c7;
    ram_cell[    1367] = 32'h0;  // 32'h201cd1e9;
    ram_cell[    1368] = 32'h0;  // 32'hc986eb2b;
    ram_cell[    1369] = 32'h0;  // 32'h9f17a61c;
    ram_cell[    1370] = 32'h0;  // 32'h366f157e;
    ram_cell[    1371] = 32'h0;  // 32'ha8e0a20c;
    ram_cell[    1372] = 32'h0;  // 32'h72fc168d;
    ram_cell[    1373] = 32'h0;  // 32'h1bc734ca;
    ram_cell[    1374] = 32'h0;  // 32'hdc938f9b;
    ram_cell[    1375] = 32'h0;  // 32'h28eff31d;
    ram_cell[    1376] = 32'h0;  // 32'h088c7ce1;
    ram_cell[    1377] = 32'h0;  // 32'he001f3dd;
    ram_cell[    1378] = 32'h0;  // 32'h4f75496e;
    ram_cell[    1379] = 32'h0;  // 32'h817a7b2a;
    ram_cell[    1380] = 32'h0;  // 32'h1cbc56d6;
    ram_cell[    1381] = 32'h0;  // 32'h85f2835f;
    ram_cell[    1382] = 32'h0;  // 32'hc7ffcb30;
    ram_cell[    1383] = 32'h0;  // 32'hc75d626d;
    ram_cell[    1384] = 32'h0;  // 32'hc96375e3;
    ram_cell[    1385] = 32'h0;  // 32'ha30c3399;
    ram_cell[    1386] = 32'h0;  // 32'hbade4e52;
    ram_cell[    1387] = 32'h0;  // 32'hc749bc6a;
    ram_cell[    1388] = 32'h0;  // 32'hdc6336c0;
    ram_cell[    1389] = 32'h0;  // 32'hef39bfea;
    ram_cell[    1390] = 32'h0;  // 32'hf7ad6f29;
    ram_cell[    1391] = 32'h0;  // 32'h8c555130;
    ram_cell[    1392] = 32'h0;  // 32'h6eea3fff;
    ram_cell[    1393] = 32'h0;  // 32'h139a5eba;
    ram_cell[    1394] = 32'h0;  // 32'h5eeefc80;
    ram_cell[    1395] = 32'h0;  // 32'h969af535;
    ram_cell[    1396] = 32'h0;  // 32'h82563a5e;
    ram_cell[    1397] = 32'h0;  // 32'hb9495b3b;
    ram_cell[    1398] = 32'h0;  // 32'he0c07316;
    ram_cell[    1399] = 32'h0;  // 32'h1e5ebaae;
    ram_cell[    1400] = 32'h0;  // 32'hee64f892;
    ram_cell[    1401] = 32'h0;  // 32'h5337890b;
    ram_cell[    1402] = 32'h0;  // 32'h9ee9edbf;
    ram_cell[    1403] = 32'h0;  // 32'hc979be3a;
    ram_cell[    1404] = 32'h0;  // 32'h07f4bcd6;
    ram_cell[    1405] = 32'h0;  // 32'hbd16d35c;
    ram_cell[    1406] = 32'h0;  // 32'h3d40cb82;
    ram_cell[    1407] = 32'h0;  // 32'h3d764e22;
    ram_cell[    1408] = 32'h0;  // 32'h41de59f6;
    ram_cell[    1409] = 32'h0;  // 32'h77296134;
    ram_cell[    1410] = 32'h0;  // 32'h11ed76f9;
    ram_cell[    1411] = 32'h0;  // 32'hd6824b68;
    ram_cell[    1412] = 32'h0;  // 32'hbe028840;
    ram_cell[    1413] = 32'h0;  // 32'hc15818df;
    ram_cell[    1414] = 32'h0;  // 32'h7ce71ef0;
    ram_cell[    1415] = 32'h0;  // 32'h8994862f;
    ram_cell[    1416] = 32'h0;  // 32'h05b409db;
    ram_cell[    1417] = 32'h0;  // 32'h9f9d21bc;
    ram_cell[    1418] = 32'h0;  // 32'hd4b9053b;
    ram_cell[    1419] = 32'h0;  // 32'h14b4cfe2;
    ram_cell[    1420] = 32'h0;  // 32'hb0d4c942;
    ram_cell[    1421] = 32'h0;  // 32'h5cdb2a52;
    ram_cell[    1422] = 32'h0;  // 32'hab849a3f;
    ram_cell[    1423] = 32'h0;  // 32'heccef157;
    ram_cell[    1424] = 32'h0;  // 32'he49bb865;
    ram_cell[    1425] = 32'h0;  // 32'h4005ba42;
    ram_cell[    1426] = 32'h0;  // 32'h07ffc465;
    ram_cell[    1427] = 32'h0;  // 32'hdfefbaa3;
    ram_cell[    1428] = 32'h0;  // 32'hce42e9d9;
    ram_cell[    1429] = 32'h0;  // 32'hf9722a81;
    ram_cell[    1430] = 32'h0;  // 32'h4f2cd37b;
    ram_cell[    1431] = 32'h0;  // 32'hf6ae5e06;
    ram_cell[    1432] = 32'h0;  // 32'h0e82a5df;
    ram_cell[    1433] = 32'h0;  // 32'h1690f683;
    ram_cell[    1434] = 32'h0;  // 32'h4e238a85;
    ram_cell[    1435] = 32'h0;  // 32'hd0176acc;
    ram_cell[    1436] = 32'h0;  // 32'h44bae984;
    ram_cell[    1437] = 32'h0;  // 32'h1b9dfa10;
    ram_cell[    1438] = 32'h0;  // 32'h631b14fc;
    ram_cell[    1439] = 32'h0;  // 32'h39985aa7;
    ram_cell[    1440] = 32'h0;  // 32'h905de7f3;
    ram_cell[    1441] = 32'h0;  // 32'h82b84e08;
    ram_cell[    1442] = 32'h0;  // 32'h22fa4506;
    ram_cell[    1443] = 32'h0;  // 32'h126f14ef;
    ram_cell[    1444] = 32'h0;  // 32'hea27cf49;
    ram_cell[    1445] = 32'h0;  // 32'h3aff2508;
    ram_cell[    1446] = 32'h0;  // 32'h888ee6a6;
    ram_cell[    1447] = 32'h0;  // 32'hf05d6038;
    ram_cell[    1448] = 32'h0;  // 32'h647e391e;
    ram_cell[    1449] = 32'h0;  // 32'h4a7bafb8;
    ram_cell[    1450] = 32'h0;  // 32'hf479c791;
    ram_cell[    1451] = 32'h0;  // 32'h8f9afe1b;
    ram_cell[    1452] = 32'h0;  // 32'h75ceaf65;
    ram_cell[    1453] = 32'h0;  // 32'h78e59601;
    ram_cell[    1454] = 32'h0;  // 32'h9247a9da;
    ram_cell[    1455] = 32'h0;  // 32'ha2820472;
    ram_cell[    1456] = 32'h0;  // 32'hd28dfba4;
    ram_cell[    1457] = 32'h0;  // 32'h9422c345;
    ram_cell[    1458] = 32'h0;  // 32'he596373e;
    ram_cell[    1459] = 32'h0;  // 32'h0a571693;
    ram_cell[    1460] = 32'h0;  // 32'h434ae3dc;
    ram_cell[    1461] = 32'h0;  // 32'h1420907e;
    ram_cell[    1462] = 32'h0;  // 32'h73721333;
    ram_cell[    1463] = 32'h0;  // 32'hc486c1a5;
    ram_cell[    1464] = 32'h0;  // 32'h298c30f3;
    ram_cell[    1465] = 32'h0;  // 32'h89e9d50e;
    ram_cell[    1466] = 32'h0;  // 32'h5327696d;
    ram_cell[    1467] = 32'h0;  // 32'h6fa1f04d;
    ram_cell[    1468] = 32'h0;  // 32'hb4e19802;
    ram_cell[    1469] = 32'h0;  // 32'h01abb4ce;
    ram_cell[    1470] = 32'h0;  // 32'h121c485e;
    ram_cell[    1471] = 32'h0;  // 32'hfbc51fc3;
    ram_cell[    1472] = 32'h0;  // 32'hc0b0621e;
    ram_cell[    1473] = 32'h0;  // 32'h7a8e1290;
    ram_cell[    1474] = 32'h0;  // 32'h4db6bd78;
    ram_cell[    1475] = 32'h0;  // 32'h40e15bed;
    ram_cell[    1476] = 32'h0;  // 32'h62bab47e;
    ram_cell[    1477] = 32'h0;  // 32'h7a6f5b74;
    ram_cell[    1478] = 32'h0;  // 32'h3881304c;
    ram_cell[    1479] = 32'h0;  // 32'h4234c107;
    ram_cell[    1480] = 32'h0;  // 32'h52cd7003;
    ram_cell[    1481] = 32'h0;  // 32'hb598a68a;
    ram_cell[    1482] = 32'h0;  // 32'hbf84b838;
    ram_cell[    1483] = 32'h0;  // 32'h294cb970;
    ram_cell[    1484] = 32'h0;  // 32'haa5330f3;
    ram_cell[    1485] = 32'h0;  // 32'haa2a70cf;
    ram_cell[    1486] = 32'h0;  // 32'hc1852685;
    ram_cell[    1487] = 32'h0;  // 32'h11c61d46;
    ram_cell[    1488] = 32'h0;  // 32'hfe718eef;
    ram_cell[    1489] = 32'h0;  // 32'h3beae2e8;
    ram_cell[    1490] = 32'h0;  // 32'h147e33c6;
    ram_cell[    1491] = 32'h0;  // 32'h16e6e6df;
    ram_cell[    1492] = 32'h0;  // 32'h05a71cd2;
    ram_cell[    1493] = 32'h0;  // 32'hd60eefb0;
    ram_cell[    1494] = 32'h0;  // 32'h66ed1d7b;
    ram_cell[    1495] = 32'h0;  // 32'h90868dc2;
    ram_cell[    1496] = 32'h0;  // 32'h7231c312;
    ram_cell[    1497] = 32'h0;  // 32'he9028af8;
    ram_cell[    1498] = 32'h0;  // 32'h1a112b46;
    ram_cell[    1499] = 32'h0;  // 32'h197583d1;
    ram_cell[    1500] = 32'h0;  // 32'h97a572b3;
    ram_cell[    1501] = 32'h0;  // 32'h41bd716e;
    ram_cell[    1502] = 32'h0;  // 32'h07f2fd83;
    ram_cell[    1503] = 32'h0;  // 32'hc8309ab7;
    ram_cell[    1504] = 32'h0;  // 32'h2e2ded51;
    ram_cell[    1505] = 32'h0;  // 32'h6dc4e827;
    ram_cell[    1506] = 32'h0;  // 32'hf1384cba;
    ram_cell[    1507] = 32'h0;  // 32'h726186f4;
    ram_cell[    1508] = 32'h0;  // 32'h89625ed9;
    ram_cell[    1509] = 32'h0;  // 32'h9afd105d;
    ram_cell[    1510] = 32'h0;  // 32'h113f8feb;
    ram_cell[    1511] = 32'h0;  // 32'hecc368c6;
    ram_cell[    1512] = 32'h0;  // 32'h06deada1;
    ram_cell[    1513] = 32'h0;  // 32'hfe213767;
    ram_cell[    1514] = 32'h0;  // 32'hb69f2691;
    ram_cell[    1515] = 32'h0;  // 32'h7bd389f9;
    ram_cell[    1516] = 32'h0;  // 32'h8bcb87b6;
    ram_cell[    1517] = 32'h0;  // 32'he4a0c7a5;
    ram_cell[    1518] = 32'h0;  // 32'h59ce8f82;
    ram_cell[    1519] = 32'h0;  // 32'hf3c11c3f;
    ram_cell[    1520] = 32'h0;  // 32'h3f6745ec;
    ram_cell[    1521] = 32'h0;  // 32'h29612ff0;
    ram_cell[    1522] = 32'h0;  // 32'h4e69e6b9;
    ram_cell[    1523] = 32'h0;  // 32'h28d9a48d;
    ram_cell[    1524] = 32'h0;  // 32'hac7c4d65;
    ram_cell[    1525] = 32'h0;  // 32'h353ef721;
    ram_cell[    1526] = 32'h0;  // 32'h25b56813;
    ram_cell[    1527] = 32'h0;  // 32'hc42e30b3;
    ram_cell[    1528] = 32'h0;  // 32'hfd2012b8;
    ram_cell[    1529] = 32'h0;  // 32'h5a77a273;
    ram_cell[    1530] = 32'h0;  // 32'h8b1eb52d;
    ram_cell[    1531] = 32'h0;  // 32'h6886189f;
    ram_cell[    1532] = 32'h0;  // 32'hf46e2e67;
    ram_cell[    1533] = 32'h0;  // 32'hc81291b4;
    ram_cell[    1534] = 32'h0;  // 32'h8471f3a5;
    ram_cell[    1535] = 32'h0;  // 32'he60c8130;
    ram_cell[    1536] = 32'h0;  // 32'h7e0ea738;
    ram_cell[    1537] = 32'h0;  // 32'hef3b90af;
    ram_cell[    1538] = 32'h0;  // 32'h90f83e26;
    ram_cell[    1539] = 32'h0;  // 32'h7eebba5e;
    ram_cell[    1540] = 32'h0;  // 32'hc4a9ea3a;
    ram_cell[    1541] = 32'h0;  // 32'h3c404319;
    ram_cell[    1542] = 32'h0;  // 32'h5a8d5357;
    ram_cell[    1543] = 32'h0;  // 32'h155e0b1a;
    ram_cell[    1544] = 32'h0;  // 32'h708d8801;
    ram_cell[    1545] = 32'h0;  // 32'h0ec8fd63;
    ram_cell[    1546] = 32'h0;  // 32'h41034927;
    ram_cell[    1547] = 32'h0;  // 32'hdad8ec23;
    ram_cell[    1548] = 32'h0;  // 32'hda995e23;
    ram_cell[    1549] = 32'h0;  // 32'h939743ef;
    ram_cell[    1550] = 32'h0;  // 32'h024c45e9;
    ram_cell[    1551] = 32'h0;  // 32'h25838354;
    ram_cell[    1552] = 32'h0;  // 32'h0d086bb0;
    ram_cell[    1553] = 32'h0;  // 32'he3f8fa47;
    ram_cell[    1554] = 32'h0;  // 32'h84c60fb0;
    ram_cell[    1555] = 32'h0;  // 32'ha18ef87f;
    ram_cell[    1556] = 32'h0;  // 32'hdb2a451e;
    ram_cell[    1557] = 32'h0;  // 32'hb861c475;
    ram_cell[    1558] = 32'h0;  // 32'h8dfd4669;
    ram_cell[    1559] = 32'h0;  // 32'hcf5fb0df;
    ram_cell[    1560] = 32'h0;  // 32'hfd6c59dd;
    ram_cell[    1561] = 32'h0;  // 32'ha8730b84;
    ram_cell[    1562] = 32'h0;  // 32'he0d9b08e;
    ram_cell[    1563] = 32'h0;  // 32'h216e594b;
    ram_cell[    1564] = 32'h0;  // 32'h4c03243c;
    ram_cell[    1565] = 32'h0;  // 32'ha1f3b4f1;
    ram_cell[    1566] = 32'h0;  // 32'hb1924979;
    ram_cell[    1567] = 32'h0;  // 32'h4301b957;
    ram_cell[    1568] = 32'h0;  // 32'hfa5e1a28;
    ram_cell[    1569] = 32'h0;  // 32'h9de4489b;
    ram_cell[    1570] = 32'h0;  // 32'h03b3be54;
    ram_cell[    1571] = 32'h0;  // 32'h7fdd1009;
    ram_cell[    1572] = 32'h0;  // 32'h804efe73;
    ram_cell[    1573] = 32'h0;  // 32'h7bd80123;
    ram_cell[    1574] = 32'h0;  // 32'h3eeb21b8;
    ram_cell[    1575] = 32'h0;  // 32'hebc589ba;
    ram_cell[    1576] = 32'h0;  // 32'h111fa612;
    ram_cell[    1577] = 32'h0;  // 32'h7ff17b7b;
    ram_cell[    1578] = 32'h0;  // 32'hd1076b0f;
    ram_cell[    1579] = 32'h0;  // 32'h2cf2fb4c;
    ram_cell[    1580] = 32'h0;  // 32'h5a42e516;
    ram_cell[    1581] = 32'h0;  // 32'h990046b3;
    ram_cell[    1582] = 32'h0;  // 32'h1ceea1ee;
    ram_cell[    1583] = 32'h0;  // 32'hf94f3d3c;
    ram_cell[    1584] = 32'h0;  // 32'h65e1f0ce;
    ram_cell[    1585] = 32'h0;  // 32'h160319a1;
    ram_cell[    1586] = 32'h0;  // 32'h916c3dbf;
    ram_cell[    1587] = 32'h0;  // 32'he56732a5;
    ram_cell[    1588] = 32'h0;  // 32'h0129e969;
    ram_cell[    1589] = 32'h0;  // 32'hc27b436f;
    ram_cell[    1590] = 32'h0;  // 32'hd5a74192;
    ram_cell[    1591] = 32'h0;  // 32'h2a53ea7e;
    ram_cell[    1592] = 32'h0;  // 32'h2d553bf8;
    ram_cell[    1593] = 32'h0;  // 32'haeaaf25b;
    ram_cell[    1594] = 32'h0;  // 32'h1b8d41b4;
    ram_cell[    1595] = 32'h0;  // 32'hceb38606;
    ram_cell[    1596] = 32'h0;  // 32'hd7230591;
    ram_cell[    1597] = 32'h0;  // 32'hcebfb6ab;
    ram_cell[    1598] = 32'h0;  // 32'h16980410;
    ram_cell[    1599] = 32'h0;  // 32'h2a8f4cf5;
    ram_cell[    1600] = 32'h0;  // 32'hd1b25baf;
    ram_cell[    1601] = 32'h0;  // 32'hb7803134;
    ram_cell[    1602] = 32'h0;  // 32'h34f7ad4c;
    ram_cell[    1603] = 32'h0;  // 32'h65e39933;
    ram_cell[    1604] = 32'h0;  // 32'hb5bac474;
    ram_cell[    1605] = 32'h0;  // 32'h4ceff987;
    ram_cell[    1606] = 32'h0;  // 32'h6f0eed30;
    ram_cell[    1607] = 32'h0;  // 32'h3043040f;
    ram_cell[    1608] = 32'h0;  // 32'h19f62e8a;
    ram_cell[    1609] = 32'h0;  // 32'hfbb6c88a;
    ram_cell[    1610] = 32'h0;  // 32'ha8a20644;
    ram_cell[    1611] = 32'h0;  // 32'h2ec3a591;
    ram_cell[    1612] = 32'h0;  // 32'h4271e76c;
    ram_cell[    1613] = 32'h0;  // 32'h3f3e65b9;
    ram_cell[    1614] = 32'h0;  // 32'hf40defec;
    ram_cell[    1615] = 32'h0;  // 32'h2d843d31;
    ram_cell[    1616] = 32'h0;  // 32'h23008e66;
    ram_cell[    1617] = 32'h0;  // 32'hcfde02ce;
    ram_cell[    1618] = 32'h0;  // 32'h53a148dc;
    ram_cell[    1619] = 32'h0;  // 32'h3577b6a4;
    ram_cell[    1620] = 32'h0;  // 32'ha709ea16;
    ram_cell[    1621] = 32'h0;  // 32'h68e8a5b5;
    ram_cell[    1622] = 32'h0;  // 32'hc016095c;
    ram_cell[    1623] = 32'h0;  // 32'h32014834;
    ram_cell[    1624] = 32'h0;  // 32'hab775be4;
    ram_cell[    1625] = 32'h0;  // 32'hb04358f0;
    ram_cell[    1626] = 32'h0;  // 32'h02861adf;
    ram_cell[    1627] = 32'h0;  // 32'h52c32ba9;
    ram_cell[    1628] = 32'h0;  // 32'h3c63688c;
    ram_cell[    1629] = 32'h0;  // 32'haf41a83e;
    ram_cell[    1630] = 32'h0;  // 32'hb4317eef;
    ram_cell[    1631] = 32'h0;  // 32'h6a0819d0;
    ram_cell[    1632] = 32'h0;  // 32'hceb07f09;
    ram_cell[    1633] = 32'h0;  // 32'h6c3993df;
    ram_cell[    1634] = 32'h0;  // 32'hb2992561;
    ram_cell[    1635] = 32'h0;  // 32'h4ef89fdb;
    ram_cell[    1636] = 32'h0;  // 32'h90f7891a;
    ram_cell[    1637] = 32'h0;  // 32'hee46b0fb;
    ram_cell[    1638] = 32'h0;  // 32'h0850f58a;
    ram_cell[    1639] = 32'h0;  // 32'h4da8573f;
    ram_cell[    1640] = 32'h0;  // 32'ha290135a;
    ram_cell[    1641] = 32'h0;  // 32'h442fdf32;
    ram_cell[    1642] = 32'h0;  // 32'h95838d14;
    ram_cell[    1643] = 32'h0;  // 32'h2dfa3122;
    ram_cell[    1644] = 32'h0;  // 32'hce5eb30d;
    ram_cell[    1645] = 32'h0;  // 32'h1c29e4bd;
    ram_cell[    1646] = 32'h0;  // 32'h8ccdd3aa;
    ram_cell[    1647] = 32'h0;  // 32'haa97fbbf;
    ram_cell[    1648] = 32'h0;  // 32'h6337005e;
    ram_cell[    1649] = 32'h0;  // 32'h95a3ab41;
    ram_cell[    1650] = 32'h0;  // 32'h58fe1e43;
    ram_cell[    1651] = 32'h0;  // 32'h8ace14f1;
    ram_cell[    1652] = 32'h0;  // 32'hb38a182a;
    ram_cell[    1653] = 32'h0;  // 32'h6ddea8a0;
    ram_cell[    1654] = 32'h0;  // 32'ha9473709;
    ram_cell[    1655] = 32'h0;  // 32'hf157a570;
    ram_cell[    1656] = 32'h0;  // 32'h9eed1e76;
    ram_cell[    1657] = 32'h0;  // 32'hda430aeb;
    ram_cell[    1658] = 32'h0;  // 32'h88cf4988;
    ram_cell[    1659] = 32'h0;  // 32'hee5431d8;
    ram_cell[    1660] = 32'h0;  // 32'h4001c3c2;
    ram_cell[    1661] = 32'h0;  // 32'h2f5cf3a7;
    ram_cell[    1662] = 32'h0;  // 32'h31e10d0c;
    ram_cell[    1663] = 32'h0;  // 32'he8c1bc78;
    ram_cell[    1664] = 32'h0;  // 32'hb3c51e95;
    ram_cell[    1665] = 32'h0;  // 32'h7a09d7f5;
    ram_cell[    1666] = 32'h0;  // 32'h236bf229;
    ram_cell[    1667] = 32'h0;  // 32'h560809b0;
    ram_cell[    1668] = 32'h0;  // 32'hb95eaa1a;
    ram_cell[    1669] = 32'h0;  // 32'h6d3af7be;
    ram_cell[    1670] = 32'h0;  // 32'h06496c9f;
    ram_cell[    1671] = 32'h0;  // 32'h519a0d32;
    ram_cell[    1672] = 32'h0;  // 32'h8ef7a9cb;
    ram_cell[    1673] = 32'h0;  // 32'h018f3a99;
    ram_cell[    1674] = 32'h0;  // 32'h9663d32a;
    ram_cell[    1675] = 32'h0;  // 32'hb1b95006;
    ram_cell[    1676] = 32'h0;  // 32'h26061414;
    ram_cell[    1677] = 32'h0;  // 32'hdecba0b5;
    ram_cell[    1678] = 32'h0;  // 32'he6740e8d;
    ram_cell[    1679] = 32'h0;  // 32'h629ab328;
    ram_cell[    1680] = 32'h0;  // 32'h4326e1da;
    ram_cell[    1681] = 32'h0;  // 32'hb80ac2c2;
    ram_cell[    1682] = 32'h0;  // 32'heaf1468a;
    ram_cell[    1683] = 32'h0;  // 32'h060e1287;
    ram_cell[    1684] = 32'h0;  // 32'heaa30193;
    ram_cell[    1685] = 32'h0;  // 32'h7e64bf51;
    ram_cell[    1686] = 32'h0;  // 32'h077fa38e;
    ram_cell[    1687] = 32'h0;  // 32'he656033f;
    ram_cell[    1688] = 32'h0;  // 32'h5ce972b1;
    ram_cell[    1689] = 32'h0;  // 32'h0fa4034c;
    ram_cell[    1690] = 32'h0;  // 32'h601ddacd;
    ram_cell[    1691] = 32'h0;  // 32'h860bb8b0;
    ram_cell[    1692] = 32'h0;  // 32'h461d6b41;
    ram_cell[    1693] = 32'h0;  // 32'h2560c92e;
    ram_cell[    1694] = 32'h0;  // 32'hdf9aa22b;
    ram_cell[    1695] = 32'h0;  // 32'hb786896f;
    ram_cell[    1696] = 32'h0;  // 32'h93fd04a9;
    ram_cell[    1697] = 32'h0;  // 32'h4208d2c6;
    ram_cell[    1698] = 32'h0;  // 32'ha152d834;
    ram_cell[    1699] = 32'h0;  // 32'ha3a4da1a;
    ram_cell[    1700] = 32'h0;  // 32'h4bef41db;
    ram_cell[    1701] = 32'h0;  // 32'ha4f1b77b;
    ram_cell[    1702] = 32'h0;  // 32'hd6bb1731;
    ram_cell[    1703] = 32'h0;  // 32'he3f9248e;
    ram_cell[    1704] = 32'h0;  // 32'h9d959028;
    ram_cell[    1705] = 32'h0;  // 32'h358f8398;
    ram_cell[    1706] = 32'h0;  // 32'h50a184bb;
    ram_cell[    1707] = 32'h0;  // 32'h447df54f;
    ram_cell[    1708] = 32'h0;  // 32'hd53624f0;
    ram_cell[    1709] = 32'h0;  // 32'h5e0d1b7d;
    ram_cell[    1710] = 32'h0;  // 32'h5c92f008;
    ram_cell[    1711] = 32'h0;  // 32'h76c3fb68;
    ram_cell[    1712] = 32'h0;  // 32'h6ab54338;
    ram_cell[    1713] = 32'h0;  // 32'h4c9d0199;
    ram_cell[    1714] = 32'h0;  // 32'h52abca77;
    ram_cell[    1715] = 32'h0;  // 32'h273627da;
    ram_cell[    1716] = 32'h0;  // 32'h8479abef;
    ram_cell[    1717] = 32'h0;  // 32'h0dff5669;
    ram_cell[    1718] = 32'h0;  // 32'h123de16c;
    ram_cell[    1719] = 32'h0;  // 32'h9dba707c;
    ram_cell[    1720] = 32'h0;  // 32'h9fa737ac;
    ram_cell[    1721] = 32'h0;  // 32'h768a9f59;
    ram_cell[    1722] = 32'h0;  // 32'h192558ae;
    ram_cell[    1723] = 32'h0;  // 32'ha2978cc0;
    ram_cell[    1724] = 32'h0;  // 32'h1b709356;
    ram_cell[    1725] = 32'h0;  // 32'hcf262610;
    ram_cell[    1726] = 32'h0;  // 32'ha1d990c5;
    ram_cell[    1727] = 32'h0;  // 32'h3534d591;
    ram_cell[    1728] = 32'h0;  // 32'h613c5839;
    ram_cell[    1729] = 32'h0;  // 32'he79d4c1e;
    ram_cell[    1730] = 32'h0;  // 32'h4845dabf;
    ram_cell[    1731] = 32'h0;  // 32'h2d88e805;
    ram_cell[    1732] = 32'h0;  // 32'h04bc3525;
    ram_cell[    1733] = 32'h0;  // 32'hf2f278b6;
    ram_cell[    1734] = 32'h0;  // 32'hd4ec704a;
    ram_cell[    1735] = 32'h0;  // 32'h7f1c829b;
    ram_cell[    1736] = 32'h0;  // 32'h68b4b6f8;
    ram_cell[    1737] = 32'h0;  // 32'h845ea9f6;
    ram_cell[    1738] = 32'h0;  // 32'h0298fe31;
    ram_cell[    1739] = 32'h0;  // 32'h9ac074e2;
    ram_cell[    1740] = 32'h0;  // 32'h3fed5390;
    ram_cell[    1741] = 32'h0;  // 32'hc65b365a;
    ram_cell[    1742] = 32'h0;  // 32'hc52e20b5;
    ram_cell[    1743] = 32'h0;  // 32'h275bddf3;
    ram_cell[    1744] = 32'h0;  // 32'h53a3f1ec;
    ram_cell[    1745] = 32'h0;  // 32'h2a2b2b03;
    ram_cell[    1746] = 32'h0;  // 32'h1de8e131;
    ram_cell[    1747] = 32'h0;  // 32'h672ad780;
    ram_cell[    1748] = 32'h0;  // 32'h3d91db26;
    ram_cell[    1749] = 32'h0;  // 32'h67e524f7;
    ram_cell[    1750] = 32'h0;  // 32'h9331c9a6;
    ram_cell[    1751] = 32'h0;  // 32'h0798878d;
    ram_cell[    1752] = 32'h0;  // 32'h6c58dbb7;
    ram_cell[    1753] = 32'h0;  // 32'h8dacb311;
    ram_cell[    1754] = 32'h0;  // 32'h09bbf5fd;
    ram_cell[    1755] = 32'h0;  // 32'h718b5e81;
    ram_cell[    1756] = 32'h0;  // 32'h770368d5;
    ram_cell[    1757] = 32'h0;  // 32'ha101a991;
    ram_cell[    1758] = 32'h0;  // 32'h371350e6;
    ram_cell[    1759] = 32'h0;  // 32'hadbc48d1;
    ram_cell[    1760] = 32'h0;  // 32'h9d62ee5e;
    ram_cell[    1761] = 32'h0;  // 32'h1f396c22;
    ram_cell[    1762] = 32'h0;  // 32'h4b1363ee;
    ram_cell[    1763] = 32'h0;  // 32'hec7a3e0b;
    ram_cell[    1764] = 32'h0;  // 32'ha8740eef;
    ram_cell[    1765] = 32'h0;  // 32'h4718aca9;
    ram_cell[    1766] = 32'h0;  // 32'ha1e31369;
    ram_cell[    1767] = 32'h0;  // 32'h2ace79f6;
    ram_cell[    1768] = 32'h0;  // 32'h96e59ab0;
    ram_cell[    1769] = 32'h0;  // 32'hf41cd081;
    ram_cell[    1770] = 32'h0;  // 32'hd6edcaea;
    ram_cell[    1771] = 32'h0;  // 32'h2ef68a41;
    ram_cell[    1772] = 32'h0;  // 32'h7ca3ef10;
    ram_cell[    1773] = 32'h0;  // 32'h0a80efdc;
    ram_cell[    1774] = 32'h0;  // 32'hf3a14ae7;
    ram_cell[    1775] = 32'h0;  // 32'h743503f5;
    ram_cell[    1776] = 32'h0;  // 32'h8eb87874;
    ram_cell[    1777] = 32'h0;  // 32'he3d0b78a;
    ram_cell[    1778] = 32'h0;  // 32'h6db5e016;
    ram_cell[    1779] = 32'h0;  // 32'h1031ca9e;
    ram_cell[    1780] = 32'h0;  // 32'h947e99ea;
    ram_cell[    1781] = 32'h0;  // 32'h2cf81ce4;
    ram_cell[    1782] = 32'h0;  // 32'h1b29d88d;
    ram_cell[    1783] = 32'h0;  // 32'h3d0239ab;
    ram_cell[    1784] = 32'h0;  // 32'hbd99e6cd;
    ram_cell[    1785] = 32'h0;  // 32'h829e6a9d;
    ram_cell[    1786] = 32'h0;  // 32'h991eab51;
    ram_cell[    1787] = 32'h0;  // 32'h954b57a0;
    ram_cell[    1788] = 32'h0;  // 32'hec5cffae;
    ram_cell[    1789] = 32'h0;  // 32'h8715130c;
    ram_cell[    1790] = 32'h0;  // 32'h77e4d863;
    ram_cell[    1791] = 32'h0;  // 32'h9a86711b;
    ram_cell[    1792] = 32'h0;  // 32'he3c28adc;
    ram_cell[    1793] = 32'h0;  // 32'h01444712;
    ram_cell[    1794] = 32'h0;  // 32'ha4b1df92;
    ram_cell[    1795] = 32'h0;  // 32'he676c6dd;
    ram_cell[    1796] = 32'h0;  // 32'h6213e8a6;
    ram_cell[    1797] = 32'h0;  // 32'h73832294;
    ram_cell[    1798] = 32'h0;  // 32'hacc104b2;
    ram_cell[    1799] = 32'h0;  // 32'hdde13454;
    ram_cell[    1800] = 32'h0;  // 32'haf61c30e;
    ram_cell[    1801] = 32'h0;  // 32'h40931223;
    ram_cell[    1802] = 32'h0;  // 32'hdad22db8;
    ram_cell[    1803] = 32'h0;  // 32'h9ceba3cf;
    ram_cell[    1804] = 32'h0;  // 32'hecc87e64;
    ram_cell[    1805] = 32'h0;  // 32'h3ea13c63;
    ram_cell[    1806] = 32'h0;  // 32'h7fa2f3bd;
    ram_cell[    1807] = 32'h0;  // 32'h1ecbd6ec;
    ram_cell[    1808] = 32'h0;  // 32'h6ed3dd2c;
    ram_cell[    1809] = 32'h0;  // 32'h2629a2ab;
    ram_cell[    1810] = 32'h0;  // 32'h0258b794;
    ram_cell[    1811] = 32'h0;  // 32'h4b4e2511;
    ram_cell[    1812] = 32'h0;  // 32'hc032a734;
    ram_cell[    1813] = 32'h0;  // 32'h6a9ea314;
    ram_cell[    1814] = 32'h0;  // 32'hf3020a38;
    ram_cell[    1815] = 32'h0;  // 32'hdd64bffd;
    ram_cell[    1816] = 32'h0;  // 32'h2de450b2;
    ram_cell[    1817] = 32'h0;  // 32'hd621a2a9;
    ram_cell[    1818] = 32'h0;  // 32'h1f663060;
    ram_cell[    1819] = 32'h0;  // 32'h98a958cb;
    ram_cell[    1820] = 32'h0;  // 32'h8f1a315c;
    ram_cell[    1821] = 32'h0;  // 32'h25dd2715;
    ram_cell[    1822] = 32'h0;  // 32'haa9fba46;
    ram_cell[    1823] = 32'h0;  // 32'hf08db45e;
    ram_cell[    1824] = 32'h0;  // 32'hd7ae5427;
    ram_cell[    1825] = 32'h0;  // 32'hddd683ae;
    ram_cell[    1826] = 32'h0;  // 32'hf805103c;
    ram_cell[    1827] = 32'h0;  // 32'hae4a31ae;
    ram_cell[    1828] = 32'h0;  // 32'h7f7d6158;
    ram_cell[    1829] = 32'h0;  // 32'h61decff4;
    ram_cell[    1830] = 32'h0;  // 32'h39d8e1b7;
    ram_cell[    1831] = 32'h0;  // 32'hc29660c2;
    ram_cell[    1832] = 32'h0;  // 32'ha44c987c;
    ram_cell[    1833] = 32'h0;  // 32'hd97e7378;
    ram_cell[    1834] = 32'h0;  // 32'h5de0a8ff;
    ram_cell[    1835] = 32'h0;  // 32'h282a6df1;
    ram_cell[    1836] = 32'h0;  // 32'hf49df4f5;
    ram_cell[    1837] = 32'h0;  // 32'h5736a364;
    ram_cell[    1838] = 32'h0;  // 32'h669b6c05;
    ram_cell[    1839] = 32'h0;  // 32'h185e377a;
    ram_cell[    1840] = 32'h0;  // 32'h10e633f6;
    ram_cell[    1841] = 32'h0;  // 32'h1873ed0c;
    ram_cell[    1842] = 32'h0;  // 32'ha94d5c0b;
    ram_cell[    1843] = 32'h0;  // 32'h4c7fac8e;
    ram_cell[    1844] = 32'h0;  // 32'hab010172;
    ram_cell[    1845] = 32'h0;  // 32'h03a1331f;
    ram_cell[    1846] = 32'h0;  // 32'h940490a5;
    ram_cell[    1847] = 32'h0;  // 32'h234c2414;
    ram_cell[    1848] = 32'h0;  // 32'h392d7075;
    ram_cell[    1849] = 32'h0;  // 32'hb0ccac54;
    ram_cell[    1850] = 32'h0;  // 32'h88090bbb;
    ram_cell[    1851] = 32'h0;  // 32'habd10354;
    ram_cell[    1852] = 32'h0;  // 32'h1d98fbe7;
    ram_cell[    1853] = 32'h0;  // 32'h1beda1bf;
    ram_cell[    1854] = 32'h0;  // 32'haf647ccc;
    ram_cell[    1855] = 32'h0;  // 32'hb9d906e7;
    ram_cell[    1856] = 32'h0;  // 32'h7c8fa04b;
    ram_cell[    1857] = 32'h0;  // 32'h2bebf4f9;
    ram_cell[    1858] = 32'h0;  // 32'hb487ebb8;
    ram_cell[    1859] = 32'h0;  // 32'h128e8ddb;
    ram_cell[    1860] = 32'h0;  // 32'h95b00dd6;
    ram_cell[    1861] = 32'h0;  // 32'h5cda460a;
    ram_cell[    1862] = 32'h0;  // 32'ha6cd8428;
    ram_cell[    1863] = 32'h0;  // 32'he9f16293;
    ram_cell[    1864] = 32'h0;  // 32'h53469cce;
    ram_cell[    1865] = 32'h0;  // 32'hc78dfd77;
    ram_cell[    1866] = 32'h0;  // 32'hdfc84783;
    ram_cell[    1867] = 32'h0;  // 32'h4164d32f;
    ram_cell[    1868] = 32'h0;  // 32'h98e31164;
    ram_cell[    1869] = 32'h0;  // 32'ha59885a9;
    ram_cell[    1870] = 32'h0;  // 32'h0ca8c64e;
    ram_cell[    1871] = 32'h0;  // 32'h7a686e39;
    ram_cell[    1872] = 32'h0;  // 32'h1e3281d4;
    ram_cell[    1873] = 32'h0;  // 32'h805d4c7a;
    ram_cell[    1874] = 32'h0;  // 32'h03af2cf2;
    ram_cell[    1875] = 32'h0;  // 32'h56f8a79b;
    ram_cell[    1876] = 32'h0;  // 32'h3e246032;
    ram_cell[    1877] = 32'h0;  // 32'h3d2f0c93;
    ram_cell[    1878] = 32'h0;  // 32'h3117a3ad;
    ram_cell[    1879] = 32'h0;  // 32'h873c7c25;
    ram_cell[    1880] = 32'h0;  // 32'hedfc74d7;
    ram_cell[    1881] = 32'h0;  // 32'ha772d1a7;
    ram_cell[    1882] = 32'h0;  // 32'ha14dd912;
    ram_cell[    1883] = 32'h0;  // 32'h31c9ece3;
    ram_cell[    1884] = 32'h0;  // 32'hdb34f3d2;
    ram_cell[    1885] = 32'h0;  // 32'h7315d5ec;
    ram_cell[    1886] = 32'h0;  // 32'ha3d6bd13;
    ram_cell[    1887] = 32'h0;  // 32'h6dfa98f4;
    ram_cell[    1888] = 32'h0;  // 32'h5da889f5;
    ram_cell[    1889] = 32'h0;  // 32'ha58291ef;
    ram_cell[    1890] = 32'h0;  // 32'he026f263;
    ram_cell[    1891] = 32'h0;  // 32'hf35ecf09;
    ram_cell[    1892] = 32'h0;  // 32'h4067d6af;
    ram_cell[    1893] = 32'h0;  // 32'heefa92ae;
    ram_cell[    1894] = 32'h0;  // 32'h3cb88c17;
    ram_cell[    1895] = 32'h0;  // 32'hc2958192;
    ram_cell[    1896] = 32'h0;  // 32'hd71a67ba;
    ram_cell[    1897] = 32'h0;  // 32'hb6913dbe;
    ram_cell[    1898] = 32'h0;  // 32'h3ee4d269;
    ram_cell[    1899] = 32'h0;  // 32'hab355c59;
    ram_cell[    1900] = 32'h0;  // 32'heab2c861;
    ram_cell[    1901] = 32'h0;  // 32'h717735c4;
    ram_cell[    1902] = 32'h0;  // 32'h929176ec;
    ram_cell[    1903] = 32'h0;  // 32'ha5f21219;
    ram_cell[    1904] = 32'h0;  // 32'hef1d27f7;
    ram_cell[    1905] = 32'h0;  // 32'hc0ec6826;
    ram_cell[    1906] = 32'h0;  // 32'h438a0e3f;
    ram_cell[    1907] = 32'h0;  // 32'h04bd76a9;
    ram_cell[    1908] = 32'h0;  // 32'h1d72eb6f;
    ram_cell[    1909] = 32'h0;  // 32'hb06d4095;
    ram_cell[    1910] = 32'h0;  // 32'h616430c0;
    ram_cell[    1911] = 32'h0;  // 32'h70ecd86f;
    ram_cell[    1912] = 32'h0;  // 32'hee3494d8;
    ram_cell[    1913] = 32'h0;  // 32'h1349c4b8;
    ram_cell[    1914] = 32'h0;  // 32'h02b109bb;
    ram_cell[    1915] = 32'h0;  // 32'h52e70e27;
    ram_cell[    1916] = 32'h0;  // 32'h2770bbfe;
    ram_cell[    1917] = 32'h0;  // 32'hc0bb4867;
    ram_cell[    1918] = 32'h0;  // 32'hf23d35e8;
    ram_cell[    1919] = 32'h0;  // 32'hfd724e2b;
    ram_cell[    1920] = 32'h0;  // 32'h0c094008;
    ram_cell[    1921] = 32'h0;  // 32'h14a1736b;
    ram_cell[    1922] = 32'h0;  // 32'h6cd4f80b;
    ram_cell[    1923] = 32'h0;  // 32'h1ac7c61f;
    ram_cell[    1924] = 32'h0;  // 32'h645c7439;
    ram_cell[    1925] = 32'h0;  // 32'hc2949e31;
    ram_cell[    1926] = 32'h0;  // 32'h5cdd915d;
    ram_cell[    1927] = 32'h0;  // 32'h5790913a;
    ram_cell[    1928] = 32'h0;  // 32'hf0e25b9c;
    ram_cell[    1929] = 32'h0;  // 32'h452d8ee4;
    ram_cell[    1930] = 32'h0;  // 32'h00fb8446;
    ram_cell[    1931] = 32'h0;  // 32'hd57f7aae;
    ram_cell[    1932] = 32'h0;  // 32'h7ce2125d;
    ram_cell[    1933] = 32'h0;  // 32'h51763e42;
    ram_cell[    1934] = 32'h0;  // 32'h79a6a54f;
    ram_cell[    1935] = 32'h0;  // 32'h1e0685ad;
    ram_cell[    1936] = 32'h0;  // 32'h50123796;
    ram_cell[    1937] = 32'h0;  // 32'hca148391;
    ram_cell[    1938] = 32'h0;  // 32'h81cabd75;
    ram_cell[    1939] = 32'h0;  // 32'h0e15cfb1;
    ram_cell[    1940] = 32'h0;  // 32'h47e3bf5e;
    ram_cell[    1941] = 32'h0;  // 32'hc1951f4b;
    ram_cell[    1942] = 32'h0;  // 32'h5f95f64e;
    ram_cell[    1943] = 32'h0;  // 32'h0ddecb48;
    ram_cell[    1944] = 32'h0;  // 32'ha973e441;
    ram_cell[    1945] = 32'h0;  // 32'hdcb2e73f;
    ram_cell[    1946] = 32'h0;  // 32'h10913440;
    ram_cell[    1947] = 32'h0;  // 32'hd8110f76;
    ram_cell[    1948] = 32'h0;  // 32'hdaec12f3;
    ram_cell[    1949] = 32'h0;  // 32'h7e2a081d;
    ram_cell[    1950] = 32'h0;  // 32'hbbdc749f;
    ram_cell[    1951] = 32'h0;  // 32'h09925be4;
    ram_cell[    1952] = 32'h0;  // 32'h602944c9;
    ram_cell[    1953] = 32'h0;  // 32'h6cd9d32e;
    ram_cell[    1954] = 32'h0;  // 32'h9a0f66a6;
    ram_cell[    1955] = 32'h0;  // 32'hc02ed524;
    ram_cell[    1956] = 32'h0;  // 32'h9f47e812;
    ram_cell[    1957] = 32'h0;  // 32'h634b7969;
    ram_cell[    1958] = 32'h0;  // 32'hc1a94404;
    ram_cell[    1959] = 32'h0;  // 32'he1260aa3;
    ram_cell[    1960] = 32'h0;  // 32'h039b25b1;
    ram_cell[    1961] = 32'h0;  // 32'h3afab491;
    ram_cell[    1962] = 32'h0;  // 32'heda094c6;
    ram_cell[    1963] = 32'h0;  // 32'ha143997d;
    ram_cell[    1964] = 32'h0;  // 32'h4fc1619f;
    ram_cell[    1965] = 32'h0;  // 32'h1801ee66;
    ram_cell[    1966] = 32'h0;  // 32'ha926ca54;
    ram_cell[    1967] = 32'h0;  // 32'h6a026fc3;
    ram_cell[    1968] = 32'h0;  // 32'he30ade59;
    ram_cell[    1969] = 32'h0;  // 32'hdd2612fa;
    ram_cell[    1970] = 32'h0;  // 32'h586f2fe9;
    ram_cell[    1971] = 32'h0;  // 32'h6a1e0181;
    ram_cell[    1972] = 32'h0;  // 32'h4a58601b;
    ram_cell[    1973] = 32'h0;  // 32'h0522e7cb;
    ram_cell[    1974] = 32'h0;  // 32'h2f14a6e0;
    ram_cell[    1975] = 32'h0;  // 32'h59cbfd60;
    ram_cell[    1976] = 32'h0;  // 32'hf5dfaed3;
    ram_cell[    1977] = 32'h0;  // 32'hcf3b1acb;
    ram_cell[    1978] = 32'h0;  // 32'hbfc0e30f;
    ram_cell[    1979] = 32'h0;  // 32'h26d7c6f7;
    ram_cell[    1980] = 32'h0;  // 32'hc5b06feb;
    ram_cell[    1981] = 32'h0;  // 32'h0bede05c;
    ram_cell[    1982] = 32'h0;  // 32'hbe9cbcd6;
    ram_cell[    1983] = 32'h0;  // 32'ha3312dc7;
    ram_cell[    1984] = 32'h0;  // 32'ha56bbd45;
    ram_cell[    1985] = 32'h0;  // 32'h05e3f093;
    ram_cell[    1986] = 32'h0;  // 32'h7c37d09c;
    ram_cell[    1987] = 32'h0;  // 32'h7c9c8fee;
    ram_cell[    1988] = 32'h0;  // 32'h36e7f76b;
    ram_cell[    1989] = 32'h0;  // 32'hde71e072;
    ram_cell[    1990] = 32'h0;  // 32'h96086858;
    ram_cell[    1991] = 32'h0;  // 32'h609da34e;
    ram_cell[    1992] = 32'h0;  // 32'hf7b157a1;
    ram_cell[    1993] = 32'h0;  // 32'h84e484d2;
    ram_cell[    1994] = 32'h0;  // 32'h09a96f4d;
    ram_cell[    1995] = 32'h0;  // 32'h80a1832b;
    ram_cell[    1996] = 32'h0;  // 32'h685e53fe;
    ram_cell[    1997] = 32'h0;  // 32'hfcd324da;
    ram_cell[    1998] = 32'h0;  // 32'hc7013352;
    ram_cell[    1999] = 32'h0;  // 32'h2f563ff4;
    ram_cell[    2000] = 32'h0;  // 32'h7b7c296a;
    ram_cell[    2001] = 32'h0;  // 32'h20dad9b8;
    ram_cell[    2002] = 32'h0;  // 32'hbaf3ad75;
    ram_cell[    2003] = 32'h0;  // 32'h59b24563;
    ram_cell[    2004] = 32'h0;  // 32'h8eae102c;
    ram_cell[    2005] = 32'h0;  // 32'h69b8e1f6;
    ram_cell[    2006] = 32'h0;  // 32'h26272d56;
    ram_cell[    2007] = 32'h0;  // 32'he2424d67;
    ram_cell[    2008] = 32'h0;  // 32'h47eb5487;
    ram_cell[    2009] = 32'h0;  // 32'h43bedb35;
    ram_cell[    2010] = 32'h0;  // 32'h0b8478dc;
    ram_cell[    2011] = 32'h0;  // 32'h3e6a6bad;
    ram_cell[    2012] = 32'h0;  // 32'hba7731fa;
    ram_cell[    2013] = 32'h0;  // 32'h62a606b5;
    ram_cell[    2014] = 32'h0;  // 32'hdb3a5f3b;
    ram_cell[    2015] = 32'h0;  // 32'h23ea1532;
    ram_cell[    2016] = 32'h0;  // 32'h4dcfb6dc;
    ram_cell[    2017] = 32'h0;  // 32'h00de77c3;
    ram_cell[    2018] = 32'h0;  // 32'hac71b9b5;
    ram_cell[    2019] = 32'h0;  // 32'h433c557c;
    ram_cell[    2020] = 32'h0;  // 32'h605cb39c;
    ram_cell[    2021] = 32'h0;  // 32'h586d92b3;
    ram_cell[    2022] = 32'h0;  // 32'hc69a0297;
    ram_cell[    2023] = 32'h0;  // 32'h420cbe2a;
    ram_cell[    2024] = 32'h0;  // 32'hb94c7037;
    ram_cell[    2025] = 32'h0;  // 32'h4ce0ce9f;
    ram_cell[    2026] = 32'h0;  // 32'ha00f84e4;
    ram_cell[    2027] = 32'h0;  // 32'h93b16e3b;
    ram_cell[    2028] = 32'h0;  // 32'h2f4309f4;
    ram_cell[    2029] = 32'h0;  // 32'h75e6bf62;
    ram_cell[    2030] = 32'h0;  // 32'hdf2233a8;
    ram_cell[    2031] = 32'h0;  // 32'hfd3960d3;
    ram_cell[    2032] = 32'h0;  // 32'h40672ca0;
    ram_cell[    2033] = 32'h0;  // 32'hbc995bc5;
    ram_cell[    2034] = 32'h0;  // 32'h7042e7cb;
    ram_cell[    2035] = 32'h0;  // 32'h77732231;
    ram_cell[    2036] = 32'h0;  // 32'h0eed8d39;
    ram_cell[    2037] = 32'h0;  // 32'h32a27765;
    ram_cell[    2038] = 32'h0;  // 32'h40ea77ca;
    ram_cell[    2039] = 32'h0;  // 32'hc8c56d2b;
    ram_cell[    2040] = 32'h0;  // 32'h76b1f940;
    ram_cell[    2041] = 32'h0;  // 32'h7901ad09;
    ram_cell[    2042] = 32'h0;  // 32'h562fbf3c;
    ram_cell[    2043] = 32'h0;  // 32'h02eb80ab;
    ram_cell[    2044] = 32'h0;  // 32'hd58b8bbe;
    ram_cell[    2045] = 32'h0;  // 32'h44713643;
    ram_cell[    2046] = 32'h0;  // 32'h2865215c;
    ram_cell[    2047] = 32'h0;  // 32'hfafbf299;
    ram_cell[    2048] = 32'h0;  // 32'hb23aa1f7;
    ram_cell[    2049] = 32'h0;  // 32'h9c4c5428;
    ram_cell[    2050] = 32'h0;  // 32'h1e1724a1;
    ram_cell[    2051] = 32'h0;  // 32'ha72d616b;
    ram_cell[    2052] = 32'h0;  // 32'h5a048482;
    ram_cell[    2053] = 32'h0;  // 32'h9fa0ee41;
    ram_cell[    2054] = 32'h0;  // 32'haba49128;
    ram_cell[    2055] = 32'h0;  // 32'hd13c4a3f;
    ram_cell[    2056] = 32'h0;  // 32'h5cfa6207;
    ram_cell[    2057] = 32'h0;  // 32'h0b999e8c;
    ram_cell[    2058] = 32'h0;  // 32'h82c29740;
    ram_cell[    2059] = 32'h0;  // 32'h4f8ba7be;
    ram_cell[    2060] = 32'h0;  // 32'h775c3c86;
    ram_cell[    2061] = 32'h0;  // 32'h10d0d8ef;
    ram_cell[    2062] = 32'h0;  // 32'h4ca85cb0;
    ram_cell[    2063] = 32'h0;  // 32'h0c3aa080;
    ram_cell[    2064] = 32'h0;  // 32'h7353efed;
    ram_cell[    2065] = 32'h0;  // 32'h4c04b69b;
    ram_cell[    2066] = 32'h0;  // 32'h6789f4cd;
    ram_cell[    2067] = 32'h0;  // 32'h35d0d9a0;
    ram_cell[    2068] = 32'h0;  // 32'hb583f4b4;
    ram_cell[    2069] = 32'h0;  // 32'h9d58afdc;
    ram_cell[    2070] = 32'h0;  // 32'h3a77258a;
    ram_cell[    2071] = 32'h0;  // 32'h780a68e1;
    ram_cell[    2072] = 32'h0;  // 32'h265aea22;
    ram_cell[    2073] = 32'h0;  // 32'hf605fbae;
    ram_cell[    2074] = 32'h0;  // 32'h9e67de77;
    ram_cell[    2075] = 32'h0;  // 32'h836fab50;
    ram_cell[    2076] = 32'h0;  // 32'hdf239d5e;
    ram_cell[    2077] = 32'h0;  // 32'h2ab8ea9e;
    ram_cell[    2078] = 32'h0;  // 32'hefdc491e;
    ram_cell[    2079] = 32'h0;  // 32'h12859842;
    ram_cell[    2080] = 32'h0;  // 32'h03cef41f;
    ram_cell[    2081] = 32'h0;  // 32'h86bfcc4e;
    ram_cell[    2082] = 32'h0;  // 32'h293646c0;
    ram_cell[    2083] = 32'h0;  // 32'hf87cacda;
    ram_cell[    2084] = 32'h0;  // 32'h5a81fbe6;
    ram_cell[    2085] = 32'h0;  // 32'h7fa5fcf9;
    ram_cell[    2086] = 32'h0;  // 32'h6c2d848e;
    ram_cell[    2087] = 32'h0;  // 32'h2062ba4f;
    ram_cell[    2088] = 32'h0;  // 32'h3625f6eb;
    ram_cell[    2089] = 32'h0;  // 32'h45abc34b;
    ram_cell[    2090] = 32'h0;  // 32'he025abef;
    ram_cell[    2091] = 32'h0;  // 32'h21d82232;
    ram_cell[    2092] = 32'h0;  // 32'h9233bdc4;
    ram_cell[    2093] = 32'h0;  // 32'hc36aa5f5;
    ram_cell[    2094] = 32'h0;  // 32'h40e379bd;
    ram_cell[    2095] = 32'h0;  // 32'h117855cf;
    ram_cell[    2096] = 32'h0;  // 32'h63df0602;
    ram_cell[    2097] = 32'h0;  // 32'h3e7ba471;
    ram_cell[    2098] = 32'h0;  // 32'hd0b26c9b;
    ram_cell[    2099] = 32'h0;  // 32'hea623246;
    ram_cell[    2100] = 32'h0;  // 32'heaecdaa7;
    ram_cell[    2101] = 32'h0;  // 32'h033b4721;
    ram_cell[    2102] = 32'h0;  // 32'hc3e01654;
    ram_cell[    2103] = 32'h0;  // 32'h2b4850f1;
    ram_cell[    2104] = 32'h0;  // 32'h94271b3c;
    ram_cell[    2105] = 32'h0;  // 32'h6664a2e7;
    ram_cell[    2106] = 32'h0;  // 32'hb9f670a0;
    ram_cell[    2107] = 32'h0;  // 32'hcf2138c0;
    ram_cell[    2108] = 32'h0;  // 32'h7ca40085;
    ram_cell[    2109] = 32'h0;  // 32'hbef57d10;
    ram_cell[    2110] = 32'h0;  // 32'hcaf3ea76;
    ram_cell[    2111] = 32'h0;  // 32'h70a09217;
    ram_cell[    2112] = 32'h0;  // 32'h8928c7b4;
    ram_cell[    2113] = 32'h0;  // 32'h4dabe9d6;
    ram_cell[    2114] = 32'h0;  // 32'hc24ff6f0;
    ram_cell[    2115] = 32'h0;  // 32'h27f795c9;
    ram_cell[    2116] = 32'h0;  // 32'h1c0e28e5;
    ram_cell[    2117] = 32'h0;  // 32'h79aebc6c;
    ram_cell[    2118] = 32'h0;  // 32'hf8fb6a1d;
    ram_cell[    2119] = 32'h0;  // 32'h139224d0;
    ram_cell[    2120] = 32'h0;  // 32'h1862ad4f;
    ram_cell[    2121] = 32'h0;  // 32'h185da6ab;
    ram_cell[    2122] = 32'h0;  // 32'h3572a602;
    ram_cell[    2123] = 32'h0;  // 32'h07f80c56;
    ram_cell[    2124] = 32'h0;  // 32'h762da69f;
    ram_cell[    2125] = 32'h0;  // 32'hd8f1298a;
    ram_cell[    2126] = 32'h0;  // 32'h05325156;
    ram_cell[    2127] = 32'h0;  // 32'he324e9e0;
    ram_cell[    2128] = 32'h0;  // 32'hc802bfd1;
    ram_cell[    2129] = 32'h0;  // 32'h9dafdc86;
    ram_cell[    2130] = 32'h0;  // 32'h24ce3dcc;
    ram_cell[    2131] = 32'h0;  // 32'hd43aaa19;
    ram_cell[    2132] = 32'h0;  // 32'hac46cfe0;
    ram_cell[    2133] = 32'h0;  // 32'hbe8f0eb8;
    ram_cell[    2134] = 32'h0;  // 32'h4834ca95;
    ram_cell[    2135] = 32'h0;  // 32'h18b39a32;
    ram_cell[    2136] = 32'h0;  // 32'h6c5975ca;
    ram_cell[    2137] = 32'h0;  // 32'h3eba0a86;
    ram_cell[    2138] = 32'h0;  // 32'h125b8568;
    ram_cell[    2139] = 32'h0;  // 32'h28eb3246;
    ram_cell[    2140] = 32'h0;  // 32'h34af3f97;
    ram_cell[    2141] = 32'h0;  // 32'hc35db62c;
    ram_cell[    2142] = 32'h0;  // 32'h087d38ca;
    ram_cell[    2143] = 32'h0;  // 32'haf495609;
    ram_cell[    2144] = 32'h0;  // 32'hc7fd6752;
    ram_cell[    2145] = 32'h0;  // 32'hc9b93020;
    ram_cell[    2146] = 32'h0;  // 32'hbf02dae7;
    ram_cell[    2147] = 32'h0;  // 32'hcaae0dac;
    ram_cell[    2148] = 32'h0;  // 32'h24556277;
    ram_cell[    2149] = 32'h0;  // 32'h19446b8c;
    ram_cell[    2150] = 32'h0;  // 32'h3c59a19b;
    ram_cell[    2151] = 32'h0;  // 32'h01242f0a;
    ram_cell[    2152] = 32'h0;  // 32'h390af4d8;
    ram_cell[    2153] = 32'h0;  // 32'ha4f28dc0;
    ram_cell[    2154] = 32'h0;  // 32'hdc12632c;
    ram_cell[    2155] = 32'h0;  // 32'h775eb217;
    ram_cell[    2156] = 32'h0;  // 32'hc4314ab6;
    ram_cell[    2157] = 32'h0;  // 32'h3855dce6;
    ram_cell[    2158] = 32'h0;  // 32'hca4e8c59;
    ram_cell[    2159] = 32'h0;  // 32'h574374b9;
    ram_cell[    2160] = 32'h0;  // 32'h428fa1b6;
    ram_cell[    2161] = 32'h0;  // 32'h0b637eaa;
    ram_cell[    2162] = 32'h0;  // 32'h86e33cd1;
    ram_cell[    2163] = 32'h0;  // 32'heb5161df;
    ram_cell[    2164] = 32'h0;  // 32'h53f22346;
    ram_cell[    2165] = 32'h0;  // 32'hd9b5640f;
    ram_cell[    2166] = 32'h0;  // 32'hff80aab8;
    ram_cell[    2167] = 32'h0;  // 32'h191c362f;
    ram_cell[    2168] = 32'h0;  // 32'h5b5af0e6;
    ram_cell[    2169] = 32'h0;  // 32'h60bf368f;
    ram_cell[    2170] = 32'h0;  // 32'h875c55fd;
    ram_cell[    2171] = 32'h0;  // 32'h88b58daa;
    ram_cell[    2172] = 32'h0;  // 32'h7dae2253;
    ram_cell[    2173] = 32'h0;  // 32'h5c967556;
    ram_cell[    2174] = 32'h0;  // 32'h3d8ed713;
    ram_cell[    2175] = 32'h0;  // 32'h7d425da8;
    ram_cell[    2176] = 32'h0;  // 32'h8343d679;
    ram_cell[    2177] = 32'h0;  // 32'h493d02f5;
    ram_cell[    2178] = 32'h0;  // 32'h84cfec09;
    ram_cell[    2179] = 32'h0;  // 32'h653209c3;
    ram_cell[    2180] = 32'h0;  // 32'h2d70d720;
    ram_cell[    2181] = 32'h0;  // 32'hbd50bc18;
    ram_cell[    2182] = 32'h0;  // 32'h64efdf41;
    ram_cell[    2183] = 32'h0;  // 32'h0ee31d41;
    ram_cell[    2184] = 32'h0;  // 32'hd052e78a;
    ram_cell[    2185] = 32'h0;  // 32'h575fb256;
    ram_cell[    2186] = 32'h0;  // 32'h89189970;
    ram_cell[    2187] = 32'h0;  // 32'hfdf10095;
    ram_cell[    2188] = 32'h0;  // 32'h89c1551e;
    ram_cell[    2189] = 32'h0;  // 32'h747aba42;
    ram_cell[    2190] = 32'h0;  // 32'h86e97383;
    ram_cell[    2191] = 32'h0;  // 32'hb9ace214;
    ram_cell[    2192] = 32'h0;  // 32'h78caaa0a;
    ram_cell[    2193] = 32'h0;  // 32'h535b438a;
    ram_cell[    2194] = 32'h0;  // 32'h774718e7;
    ram_cell[    2195] = 32'h0;  // 32'hd2b15c12;
    ram_cell[    2196] = 32'h0;  // 32'h0291dd77;
    ram_cell[    2197] = 32'h0;  // 32'he84e0507;
    ram_cell[    2198] = 32'h0;  // 32'h0b25c974;
    ram_cell[    2199] = 32'h0;  // 32'h82281e66;
    ram_cell[    2200] = 32'h0;  // 32'hc5190d1c;
    ram_cell[    2201] = 32'h0;  // 32'h43d0abbd;
    ram_cell[    2202] = 32'h0;  // 32'hf76bca0a;
    ram_cell[    2203] = 32'h0;  // 32'h1161f611;
    ram_cell[    2204] = 32'h0;  // 32'h446a9304;
    ram_cell[    2205] = 32'h0;  // 32'h40b2414a;
    ram_cell[    2206] = 32'h0;  // 32'he1c8e967;
    ram_cell[    2207] = 32'h0;  // 32'hb923088f;
    ram_cell[    2208] = 32'h0;  // 32'h71050fab;
    ram_cell[    2209] = 32'h0;  // 32'hb41f5a20;
    ram_cell[    2210] = 32'h0;  // 32'hef7ad60e;
    ram_cell[    2211] = 32'h0;  // 32'hcbe39de5;
    ram_cell[    2212] = 32'h0;  // 32'he97a904a;
    ram_cell[    2213] = 32'h0;  // 32'h89c3752e;
    ram_cell[    2214] = 32'h0;  // 32'hb2228e6e;
    ram_cell[    2215] = 32'h0;  // 32'he6a0cba4;
    ram_cell[    2216] = 32'h0;  // 32'h99af9c59;
    ram_cell[    2217] = 32'h0;  // 32'hfa3152b3;
    ram_cell[    2218] = 32'h0;  // 32'h82a76a99;
    ram_cell[    2219] = 32'h0;  // 32'h8f77ace1;
    ram_cell[    2220] = 32'h0;  // 32'h70c37aef;
    ram_cell[    2221] = 32'h0;  // 32'h9cc22c67;
    ram_cell[    2222] = 32'h0;  // 32'h32689ef8;
    ram_cell[    2223] = 32'h0;  // 32'h33ab8786;
    ram_cell[    2224] = 32'h0;  // 32'h8eb0768e;
    ram_cell[    2225] = 32'h0;  // 32'hb3cd2c42;
    ram_cell[    2226] = 32'h0;  // 32'he4bf70de;
    ram_cell[    2227] = 32'h0;  // 32'h8e2839bf;
    ram_cell[    2228] = 32'h0;  // 32'ha8767a2b;
    ram_cell[    2229] = 32'h0;  // 32'h79536434;
    ram_cell[    2230] = 32'h0;  // 32'h404e8697;
    ram_cell[    2231] = 32'h0;  // 32'h36f7357c;
    ram_cell[    2232] = 32'h0;  // 32'h2c810b31;
    ram_cell[    2233] = 32'h0;  // 32'he21aa971;
    ram_cell[    2234] = 32'h0;  // 32'ha016eed8;
    ram_cell[    2235] = 32'h0;  // 32'h52e06808;
    ram_cell[    2236] = 32'h0;  // 32'hada1f290;
    ram_cell[    2237] = 32'h0;  // 32'haa663a63;
    ram_cell[    2238] = 32'h0;  // 32'hf5366c52;
    ram_cell[    2239] = 32'h0;  // 32'hc0218d71;
    ram_cell[    2240] = 32'h0;  // 32'h89a83011;
    ram_cell[    2241] = 32'h0;  // 32'h09009234;
    ram_cell[    2242] = 32'h0;  // 32'hff5e5007;
    ram_cell[    2243] = 32'h0;  // 32'hcf72b124;
    ram_cell[    2244] = 32'h0;  // 32'h43442e45;
    ram_cell[    2245] = 32'h0;  // 32'h03978c3d;
    ram_cell[    2246] = 32'h0;  // 32'h808974c0;
    ram_cell[    2247] = 32'h0;  // 32'h41ef0686;
    ram_cell[    2248] = 32'h0;  // 32'h2fe3380f;
    ram_cell[    2249] = 32'h0;  // 32'h740bdaab;
    ram_cell[    2250] = 32'h0;  // 32'h86152491;
    ram_cell[    2251] = 32'h0;  // 32'h4aff8398;
    ram_cell[    2252] = 32'h0;  // 32'he7416c4c;
    ram_cell[    2253] = 32'h0;  // 32'h00096fb5;
    ram_cell[    2254] = 32'h0;  // 32'hfdc4138b;
    ram_cell[    2255] = 32'h0;  // 32'h9812b9b4;
    ram_cell[    2256] = 32'h0;  // 32'had2ea3d4;
    ram_cell[    2257] = 32'h0;  // 32'h51b31ca0;
    ram_cell[    2258] = 32'h0;  // 32'h44142db2;
    ram_cell[    2259] = 32'h0;  // 32'h03376b27;
    ram_cell[    2260] = 32'h0;  // 32'h22e89dcd;
    ram_cell[    2261] = 32'h0;  // 32'hef962561;
    ram_cell[    2262] = 32'h0;  // 32'hbf4438bf;
    ram_cell[    2263] = 32'h0;  // 32'h95aec07c;
    ram_cell[    2264] = 32'h0;  // 32'hca680a4e;
    ram_cell[    2265] = 32'h0;  // 32'hdc86026d;
    ram_cell[    2266] = 32'h0;  // 32'h3d854d57;
    ram_cell[    2267] = 32'h0;  // 32'h13424a3a;
    ram_cell[    2268] = 32'h0;  // 32'hc8870065;
    ram_cell[    2269] = 32'h0;  // 32'h4d622712;
    ram_cell[    2270] = 32'h0;  // 32'h628a4f60;
    ram_cell[    2271] = 32'h0;  // 32'ha9508dff;
    ram_cell[    2272] = 32'h0;  // 32'he44661c6;
    ram_cell[    2273] = 32'h0;  // 32'hc7f4ae3f;
    ram_cell[    2274] = 32'h0;  // 32'h2ebe4126;
    ram_cell[    2275] = 32'h0;  // 32'h3a309e16;
    ram_cell[    2276] = 32'h0;  // 32'hdcdd0ca5;
    ram_cell[    2277] = 32'h0;  // 32'h90f6d6da;
    ram_cell[    2278] = 32'h0;  // 32'h77d93974;
    ram_cell[    2279] = 32'h0;  // 32'h20b512b4;
    ram_cell[    2280] = 32'h0;  // 32'h723f34cb;
    ram_cell[    2281] = 32'h0;  // 32'h9bee744e;
    ram_cell[    2282] = 32'h0;  // 32'h7e24b8ed;
    ram_cell[    2283] = 32'h0;  // 32'hc4a3dc00;
    ram_cell[    2284] = 32'h0;  // 32'hb39fcebe;
    ram_cell[    2285] = 32'h0;  // 32'h2c59dc99;
    ram_cell[    2286] = 32'h0;  // 32'h3f7a9958;
    ram_cell[    2287] = 32'h0;  // 32'h8ce3074c;
    ram_cell[    2288] = 32'h0;  // 32'h034b072b;
    ram_cell[    2289] = 32'h0;  // 32'hc42fe864;
    ram_cell[    2290] = 32'h0;  // 32'hbbefde91;
    ram_cell[    2291] = 32'h0;  // 32'h1f61948f;
    ram_cell[    2292] = 32'h0;  // 32'h6ddbe530;
    ram_cell[    2293] = 32'h0;  // 32'hbbf6c705;
    ram_cell[    2294] = 32'h0;  // 32'hf10a0d27;
    ram_cell[    2295] = 32'h0;  // 32'hc0072bf9;
    ram_cell[    2296] = 32'h0;  // 32'h4ff1e3f4;
    ram_cell[    2297] = 32'h0;  // 32'h51d9f97e;
    ram_cell[    2298] = 32'h0;  // 32'h81899542;
    ram_cell[    2299] = 32'h0;  // 32'h9e1415a2;
    ram_cell[    2300] = 32'h0;  // 32'hdf0ee464;
    ram_cell[    2301] = 32'h0;  // 32'h2a5736f5;
    ram_cell[    2302] = 32'h0;  // 32'h7b18f2e5;
    ram_cell[    2303] = 32'h0;  // 32'ha795acd3;
    ram_cell[    2304] = 32'h0;  // 32'hcf66dc6d;
    ram_cell[    2305] = 32'h0;  // 32'he8727c9e;
    ram_cell[    2306] = 32'h0;  // 32'h8f6b7188;
    ram_cell[    2307] = 32'h0;  // 32'hc1bb3873;
    ram_cell[    2308] = 32'h0;  // 32'h5fe0561a;
    ram_cell[    2309] = 32'h0;  // 32'h2c368989;
    ram_cell[    2310] = 32'h0;  // 32'h03f19a97;
    ram_cell[    2311] = 32'h0;  // 32'hbc80b75c;
    ram_cell[    2312] = 32'h0;  // 32'h03f38853;
    ram_cell[    2313] = 32'h0;  // 32'ha26192a8;
    ram_cell[    2314] = 32'h0;  // 32'hac4f3937;
    ram_cell[    2315] = 32'h0;  // 32'hc46d31e6;
    ram_cell[    2316] = 32'h0;  // 32'h18e786d1;
    ram_cell[    2317] = 32'h0;  // 32'h563bc198;
    ram_cell[    2318] = 32'h0;  // 32'h50061114;
    ram_cell[    2319] = 32'h0;  // 32'hefef3382;
    ram_cell[    2320] = 32'h0;  // 32'ha0f0bc12;
    ram_cell[    2321] = 32'h0;  // 32'h6e36863f;
    ram_cell[    2322] = 32'h0;  // 32'he501c6d8;
    ram_cell[    2323] = 32'h0;  // 32'h425e45e6;
    ram_cell[    2324] = 32'h0;  // 32'hcc7dd61b;
    ram_cell[    2325] = 32'h0;  // 32'h925d7633;
    ram_cell[    2326] = 32'h0;  // 32'h22c8dd76;
    ram_cell[    2327] = 32'h0;  // 32'haa43ac9c;
    ram_cell[    2328] = 32'h0;  // 32'h1f068126;
    ram_cell[    2329] = 32'h0;  // 32'hb50c7c8f;
    ram_cell[    2330] = 32'h0;  // 32'h24444d2d;
    ram_cell[    2331] = 32'h0;  // 32'h17ceca97;
    ram_cell[    2332] = 32'h0;  // 32'h13503a3a;
    ram_cell[    2333] = 32'h0;  // 32'h21fc1d79;
    ram_cell[    2334] = 32'h0;  // 32'he5b9effd;
    ram_cell[    2335] = 32'h0;  // 32'h470018bc;
    ram_cell[    2336] = 32'h0;  // 32'h10e0c2e3;
    ram_cell[    2337] = 32'h0;  // 32'h4c36ca02;
    ram_cell[    2338] = 32'h0;  // 32'h5a544afc;
    ram_cell[    2339] = 32'h0;  // 32'h1a8cce75;
    ram_cell[    2340] = 32'h0;  // 32'hd416d17d;
    ram_cell[    2341] = 32'h0;  // 32'h498f631d;
    ram_cell[    2342] = 32'h0;  // 32'h02fd8f87;
    ram_cell[    2343] = 32'h0;  // 32'h1241bbaa;
    ram_cell[    2344] = 32'h0;  // 32'h78774e81;
    ram_cell[    2345] = 32'h0;  // 32'h9844839b;
    ram_cell[    2346] = 32'h0;  // 32'hce12d19d;
    ram_cell[    2347] = 32'h0;  // 32'hef4066af;
    ram_cell[    2348] = 32'h0;  // 32'hf457e78c;
    ram_cell[    2349] = 32'h0;  // 32'h473ea268;
    ram_cell[    2350] = 32'h0;  // 32'hd21b13b2;
    ram_cell[    2351] = 32'h0;  // 32'h094ed7b0;
    ram_cell[    2352] = 32'h0;  // 32'h3dae9bef;
    ram_cell[    2353] = 32'h0;  // 32'hc18ede7f;
    ram_cell[    2354] = 32'h0;  // 32'hfcb0c28f;
    ram_cell[    2355] = 32'h0;  // 32'hd662e81e;
    ram_cell[    2356] = 32'h0;  // 32'h2e9e122a;
    ram_cell[    2357] = 32'h0;  // 32'h98bbece3;
    ram_cell[    2358] = 32'h0;  // 32'h09c6e398;
    ram_cell[    2359] = 32'h0;  // 32'h31fa6bb6;
    ram_cell[    2360] = 32'h0;  // 32'hc01a7f37;
    ram_cell[    2361] = 32'h0;  // 32'hcd9b05c2;
    ram_cell[    2362] = 32'h0;  // 32'h7a3fad23;
    ram_cell[    2363] = 32'h0;  // 32'h1aa3cf66;
    ram_cell[    2364] = 32'h0;  // 32'h87a94542;
    ram_cell[    2365] = 32'h0;  // 32'h08fa5bbc;
    ram_cell[    2366] = 32'h0;  // 32'hba33e346;
    ram_cell[    2367] = 32'h0;  // 32'h93891a54;
    ram_cell[    2368] = 32'h0;  // 32'h306145b4;
    ram_cell[    2369] = 32'h0;  // 32'h56fa7dab;
    ram_cell[    2370] = 32'h0;  // 32'h8aa7f09b;
    ram_cell[    2371] = 32'h0;  // 32'h5f434693;
    ram_cell[    2372] = 32'h0;  // 32'h02d033b1;
    ram_cell[    2373] = 32'h0;  // 32'h3ab899e7;
    ram_cell[    2374] = 32'h0;  // 32'hacf85c9d;
    ram_cell[    2375] = 32'h0;  // 32'h4f5580ff;
    ram_cell[    2376] = 32'h0;  // 32'habcea15a;
    ram_cell[    2377] = 32'h0;  // 32'h7455b995;
    ram_cell[    2378] = 32'h0;  // 32'hdee08fae;
    ram_cell[    2379] = 32'h0;  // 32'h0431155e;
    ram_cell[    2380] = 32'h0;  // 32'h2ed07709;
    ram_cell[    2381] = 32'h0;  // 32'h16e399ae;
    ram_cell[    2382] = 32'h0;  // 32'hdfcaffa4;
    ram_cell[    2383] = 32'h0;  // 32'h2b90de61;
    ram_cell[    2384] = 32'h0;  // 32'hee8211e8;
    ram_cell[    2385] = 32'h0;  // 32'hbd1a1964;
    ram_cell[    2386] = 32'h0;  // 32'hba546297;
    ram_cell[    2387] = 32'h0;  // 32'h29634a5b;
    ram_cell[    2388] = 32'h0;  // 32'he26cf76f;
    ram_cell[    2389] = 32'h0;  // 32'h60ede301;
    ram_cell[    2390] = 32'h0;  // 32'ha9f64209;
    ram_cell[    2391] = 32'h0;  // 32'h58f731fa;
    ram_cell[    2392] = 32'h0;  // 32'hbb39a871;
    ram_cell[    2393] = 32'h0;  // 32'h31380858;
    ram_cell[    2394] = 32'h0;  // 32'h63498533;
    ram_cell[    2395] = 32'h0;  // 32'heafe8906;
    ram_cell[    2396] = 32'h0;  // 32'he987389e;
    ram_cell[    2397] = 32'h0;  // 32'hb5860513;
    ram_cell[    2398] = 32'h0;  // 32'h1eb66891;
    ram_cell[    2399] = 32'h0;  // 32'h3d495796;
    ram_cell[    2400] = 32'h0;  // 32'h14d9009c;
    ram_cell[    2401] = 32'h0;  // 32'h642cba83;
    ram_cell[    2402] = 32'h0;  // 32'h7563a988;
    ram_cell[    2403] = 32'h0;  // 32'h2837ae06;
    ram_cell[    2404] = 32'h0;  // 32'haa588ddb;
    ram_cell[    2405] = 32'h0;  // 32'h790c5954;
    ram_cell[    2406] = 32'h0;  // 32'hd978326f;
    ram_cell[    2407] = 32'h0;  // 32'h916eb6e8;
    ram_cell[    2408] = 32'h0;  // 32'hf3b7d1d2;
    ram_cell[    2409] = 32'h0;  // 32'hb5ba1eab;
    ram_cell[    2410] = 32'h0;  // 32'hf4d099f9;
    ram_cell[    2411] = 32'h0;  // 32'h23a72d3d;
    ram_cell[    2412] = 32'h0;  // 32'h04367c93;
    ram_cell[    2413] = 32'h0;  // 32'hcc3a78ff;
    ram_cell[    2414] = 32'h0;  // 32'h18f945d9;
    ram_cell[    2415] = 32'h0;  // 32'h3f393d7d;
    ram_cell[    2416] = 32'h0;  // 32'h1ed290f5;
    ram_cell[    2417] = 32'h0;  // 32'hfb18fd79;
    ram_cell[    2418] = 32'h0;  // 32'heb2aff96;
    ram_cell[    2419] = 32'h0;  // 32'he0b5f981;
    ram_cell[    2420] = 32'h0;  // 32'hf362e0c3;
    ram_cell[    2421] = 32'h0;  // 32'hd7cc7e27;
    ram_cell[    2422] = 32'h0;  // 32'h1cfcdc15;
    ram_cell[    2423] = 32'h0;  // 32'hadc5cf7a;
    ram_cell[    2424] = 32'h0;  // 32'h77d38252;
    ram_cell[    2425] = 32'h0;  // 32'h7bf83c8d;
    ram_cell[    2426] = 32'h0;  // 32'h519652b0;
    ram_cell[    2427] = 32'h0;  // 32'he39b8463;
    ram_cell[    2428] = 32'h0;  // 32'h84a910b3;
    ram_cell[    2429] = 32'h0;  // 32'h2149da12;
    ram_cell[    2430] = 32'h0;  // 32'h87de9992;
    ram_cell[    2431] = 32'h0;  // 32'h07db94db;
    ram_cell[    2432] = 32'h0;  // 32'hf5024259;
    ram_cell[    2433] = 32'h0;  // 32'ha18c177f;
    ram_cell[    2434] = 32'h0;  // 32'h23309694;
    ram_cell[    2435] = 32'h0;  // 32'h36044e43;
    ram_cell[    2436] = 32'h0;  // 32'hd00a1904;
    ram_cell[    2437] = 32'h0;  // 32'hc1914315;
    ram_cell[    2438] = 32'h0;  // 32'h2a5263de;
    ram_cell[    2439] = 32'h0;  // 32'h5450b65f;
    ram_cell[    2440] = 32'h0;  // 32'h39c6ca66;
    ram_cell[    2441] = 32'h0;  // 32'h0b32bf88;
    ram_cell[    2442] = 32'h0;  // 32'hd612a287;
    ram_cell[    2443] = 32'h0;  // 32'h6781c8db;
    ram_cell[    2444] = 32'h0;  // 32'hce1aec19;
    ram_cell[    2445] = 32'h0;  // 32'hb61fb511;
    ram_cell[    2446] = 32'h0;  // 32'hbc10c7ee;
    ram_cell[    2447] = 32'h0;  // 32'haaa1da4d;
    ram_cell[    2448] = 32'h0;  // 32'h319c0df2;
    ram_cell[    2449] = 32'h0;  // 32'h84bf457f;
    ram_cell[    2450] = 32'h0;  // 32'h33cec447;
    ram_cell[    2451] = 32'h0;  // 32'ha00e2973;
    ram_cell[    2452] = 32'h0;  // 32'h68a9b951;
    ram_cell[    2453] = 32'h0;  // 32'hb0e63756;
    ram_cell[    2454] = 32'h0;  // 32'h850977b9;
    ram_cell[    2455] = 32'h0;  // 32'ha9d1c1fd;
    ram_cell[    2456] = 32'h0;  // 32'h0bcb658a;
    ram_cell[    2457] = 32'h0;  // 32'h35c2eb27;
    ram_cell[    2458] = 32'h0;  // 32'ha6a17dae;
    ram_cell[    2459] = 32'h0;  // 32'h4f79a9a5;
    ram_cell[    2460] = 32'h0;  // 32'ha0e6abc2;
    ram_cell[    2461] = 32'h0;  // 32'h541cec9e;
    ram_cell[    2462] = 32'h0;  // 32'h181c7c5b;
    ram_cell[    2463] = 32'h0;  // 32'h5a63756b;
    ram_cell[    2464] = 32'h0;  // 32'h20ad13e4;
    ram_cell[    2465] = 32'h0;  // 32'h02d777fd;
    ram_cell[    2466] = 32'h0;  // 32'hbc362cee;
    ram_cell[    2467] = 32'h0;  // 32'h66b694f1;
    ram_cell[    2468] = 32'h0;  // 32'h02ede9d5;
    ram_cell[    2469] = 32'h0;  // 32'hca7c8604;
    ram_cell[    2470] = 32'h0;  // 32'ha22121e0;
    ram_cell[    2471] = 32'h0;  // 32'h6a237915;
    ram_cell[    2472] = 32'h0;  // 32'h8b85079e;
    ram_cell[    2473] = 32'h0;  // 32'hf07ac667;
    ram_cell[    2474] = 32'h0;  // 32'hb38f15f3;
    ram_cell[    2475] = 32'h0;  // 32'heb6dcfb5;
    ram_cell[    2476] = 32'h0;  // 32'h05f57208;
    ram_cell[    2477] = 32'h0;  // 32'he4f8a6ca;
    ram_cell[    2478] = 32'h0;  // 32'h71422beb;
    ram_cell[    2479] = 32'h0;  // 32'h11787134;
    ram_cell[    2480] = 32'h0;  // 32'h4d12a964;
    ram_cell[    2481] = 32'h0;  // 32'h3d991dc5;
    ram_cell[    2482] = 32'h0;  // 32'h53a81874;
    ram_cell[    2483] = 32'h0;  // 32'hdb897905;
    ram_cell[    2484] = 32'h0;  // 32'hc80f3bbc;
    ram_cell[    2485] = 32'h0;  // 32'hb203ab5b;
    ram_cell[    2486] = 32'h0;  // 32'h2533cc79;
    ram_cell[    2487] = 32'h0;  // 32'h2c918441;
    ram_cell[    2488] = 32'h0;  // 32'hf9950db7;
    ram_cell[    2489] = 32'h0;  // 32'ha5553224;
    ram_cell[    2490] = 32'h0;  // 32'h163931b3;
    ram_cell[    2491] = 32'h0;  // 32'hd9639ffd;
    ram_cell[    2492] = 32'h0;  // 32'h3ffbfa25;
    ram_cell[    2493] = 32'h0;  // 32'h2bfc3818;
    ram_cell[    2494] = 32'h0;  // 32'h4c649f21;
    ram_cell[    2495] = 32'h0;  // 32'h45baa9dd;
    ram_cell[    2496] = 32'h0;  // 32'h9662dd1c;
    ram_cell[    2497] = 32'h0;  // 32'h71f76667;
    ram_cell[    2498] = 32'h0;  // 32'h4d2027d6;
    ram_cell[    2499] = 32'h0;  // 32'ha9dc0ef7;
    ram_cell[    2500] = 32'h0;  // 32'h40590e01;
    ram_cell[    2501] = 32'h0;  // 32'haac764e1;
    ram_cell[    2502] = 32'h0;  // 32'h985f3e5a;
    ram_cell[    2503] = 32'h0;  // 32'hd74e1d0a;
    ram_cell[    2504] = 32'h0;  // 32'hf38e1c76;
    ram_cell[    2505] = 32'h0;  // 32'h90ed68d9;
    ram_cell[    2506] = 32'h0;  // 32'h87349f37;
    ram_cell[    2507] = 32'h0;  // 32'hd04a0e00;
    ram_cell[    2508] = 32'h0;  // 32'h93c4d1d9;
    ram_cell[    2509] = 32'h0;  // 32'h5a797f37;
    ram_cell[    2510] = 32'h0;  // 32'hc724e4f6;
    ram_cell[    2511] = 32'h0;  // 32'h202686e5;
    ram_cell[    2512] = 32'h0;  // 32'h90c27e6e;
    ram_cell[    2513] = 32'h0;  // 32'hb64291d9;
    ram_cell[    2514] = 32'h0;  // 32'h4e2f787e;
    ram_cell[    2515] = 32'h0;  // 32'h3279725f;
    ram_cell[    2516] = 32'h0;  // 32'h2e169dce;
    ram_cell[    2517] = 32'h0;  // 32'h07f6dc95;
    ram_cell[    2518] = 32'h0;  // 32'h9cb6f2af;
    ram_cell[    2519] = 32'h0;  // 32'h061dd9b6;
    ram_cell[    2520] = 32'h0;  // 32'h12ffa5e7;
    ram_cell[    2521] = 32'h0;  // 32'h9a69491a;
    ram_cell[    2522] = 32'h0;  // 32'h2ce8301c;
    ram_cell[    2523] = 32'h0;  // 32'h72922f20;
    ram_cell[    2524] = 32'h0;  // 32'h66093aaf;
    ram_cell[    2525] = 32'h0;  // 32'hedfcce59;
    ram_cell[    2526] = 32'h0;  // 32'hb3bfe3df;
    ram_cell[    2527] = 32'h0;  // 32'h7bcc3c14;
    ram_cell[    2528] = 32'h0;  // 32'h758f57ee;
    ram_cell[    2529] = 32'h0;  // 32'h0c97cd73;
    ram_cell[    2530] = 32'h0;  // 32'h44c62a54;
    ram_cell[    2531] = 32'h0;  // 32'h38aa16d6;
    ram_cell[    2532] = 32'h0;  // 32'hce29547b;
    ram_cell[    2533] = 32'h0;  // 32'h88935ce8;
    ram_cell[    2534] = 32'h0;  // 32'h95518ae4;
    ram_cell[    2535] = 32'h0;  // 32'h59b83e6f;
    ram_cell[    2536] = 32'h0;  // 32'hbb83d0f0;
    ram_cell[    2537] = 32'h0;  // 32'h3fd5d317;
    ram_cell[    2538] = 32'h0;  // 32'h5d3453e1;
    ram_cell[    2539] = 32'h0;  // 32'hefec2f3c;
    ram_cell[    2540] = 32'h0;  // 32'h42cc021f;
    ram_cell[    2541] = 32'h0;  // 32'hbf336272;
    ram_cell[    2542] = 32'h0;  // 32'h6f72df28;
    ram_cell[    2543] = 32'h0;  // 32'he35fcd42;
    ram_cell[    2544] = 32'h0;  // 32'h49816645;
    ram_cell[    2545] = 32'h0;  // 32'h7860da41;
    ram_cell[    2546] = 32'h0;  // 32'h23748327;
    ram_cell[    2547] = 32'h0;  // 32'h5d198a6c;
    ram_cell[    2548] = 32'h0;  // 32'h41f85a18;
    ram_cell[    2549] = 32'h0;  // 32'h4a095910;
    ram_cell[    2550] = 32'h0;  // 32'hc344f897;
    ram_cell[    2551] = 32'h0;  // 32'h2c751d0f;
    ram_cell[    2552] = 32'h0;  // 32'h48643c84;
    ram_cell[    2553] = 32'h0;  // 32'he615d1b3;
    ram_cell[    2554] = 32'h0;  // 32'h505194e3;
    ram_cell[    2555] = 32'h0;  // 32'h85283592;
    ram_cell[    2556] = 32'h0;  // 32'h95d37dcf;
    ram_cell[    2557] = 32'h0;  // 32'h93056f30;
    ram_cell[    2558] = 32'h0;  // 32'h700908c4;
    ram_cell[    2559] = 32'h0;  // 32'h53debc56;
    ram_cell[    2560] = 32'h0;  // 32'h07ddae70;
    ram_cell[    2561] = 32'h0;  // 32'h995aed17;
    ram_cell[    2562] = 32'h0;  // 32'h294ca739;
    ram_cell[    2563] = 32'h0;  // 32'hd61374d7;
    ram_cell[    2564] = 32'h0;  // 32'h09b2f380;
    ram_cell[    2565] = 32'h0;  // 32'h817c20ec;
    ram_cell[    2566] = 32'h0;  // 32'h50cad952;
    ram_cell[    2567] = 32'h0;  // 32'h5ba19bb2;
    ram_cell[    2568] = 32'h0;  // 32'h17438190;
    ram_cell[    2569] = 32'h0;  // 32'he654ff9e;
    ram_cell[    2570] = 32'h0;  // 32'hdc634cc8;
    ram_cell[    2571] = 32'h0;  // 32'h0eecb249;
    ram_cell[    2572] = 32'h0;  // 32'hf0a4baa0;
    ram_cell[    2573] = 32'h0;  // 32'hefd4b3f1;
    ram_cell[    2574] = 32'h0;  // 32'h221bb2b2;
    ram_cell[    2575] = 32'h0;  // 32'h7c9ec66f;
    ram_cell[    2576] = 32'h0;  // 32'hf5b6c669;
    ram_cell[    2577] = 32'h0;  // 32'h62eebf05;
    ram_cell[    2578] = 32'h0;  // 32'h1a58eb0a;
    ram_cell[    2579] = 32'h0;  // 32'h20e7f341;
    ram_cell[    2580] = 32'h0;  // 32'h56cf67a4;
    ram_cell[    2581] = 32'h0;  // 32'hce7732ac;
    ram_cell[    2582] = 32'h0;  // 32'h3ca4f237;
    ram_cell[    2583] = 32'h0;  // 32'hcd11b31b;
    ram_cell[    2584] = 32'h0;  // 32'h3d7f64a3;
    ram_cell[    2585] = 32'h0;  // 32'h6b5f7ef8;
    ram_cell[    2586] = 32'h0;  // 32'h0587a87b;
    ram_cell[    2587] = 32'h0;  // 32'hddcf5027;
    ram_cell[    2588] = 32'h0;  // 32'h61778722;
    ram_cell[    2589] = 32'h0;  // 32'h2c19a845;
    ram_cell[    2590] = 32'h0;  // 32'h783db687;
    ram_cell[    2591] = 32'h0;  // 32'h3e560cf8;
    ram_cell[    2592] = 32'h0;  // 32'hdd9a094f;
    ram_cell[    2593] = 32'h0;  // 32'h580496ca;
    ram_cell[    2594] = 32'h0;  // 32'h969ecd29;
    ram_cell[    2595] = 32'h0;  // 32'h1553f4b6;
    ram_cell[    2596] = 32'h0;  // 32'h121cd21b;
    ram_cell[    2597] = 32'h0;  // 32'h9fa99ac0;
    ram_cell[    2598] = 32'h0;  // 32'hfa43e93e;
    ram_cell[    2599] = 32'h0;  // 32'h035a44ec;
    ram_cell[    2600] = 32'h0;  // 32'hf77134b8;
    ram_cell[    2601] = 32'h0;  // 32'h5cd98552;
    ram_cell[    2602] = 32'h0;  // 32'h98f74e8d;
    ram_cell[    2603] = 32'h0;  // 32'h266da1a5;
    ram_cell[    2604] = 32'h0;  // 32'h77e03bc9;
    ram_cell[    2605] = 32'h0;  // 32'h824b3775;
    ram_cell[    2606] = 32'h0;  // 32'h9a2580e0;
    ram_cell[    2607] = 32'h0;  // 32'h1f2a8127;
    ram_cell[    2608] = 32'h0;  // 32'h38e83fc8;
    ram_cell[    2609] = 32'h0;  // 32'h04103da6;
    ram_cell[    2610] = 32'h0;  // 32'he3fbdc93;
    ram_cell[    2611] = 32'h0;  // 32'hf69f8e35;
    ram_cell[    2612] = 32'h0;  // 32'hfec4493f;
    ram_cell[    2613] = 32'h0;  // 32'h21561477;
    ram_cell[    2614] = 32'h0;  // 32'h4487c3d6;
    ram_cell[    2615] = 32'h0;  // 32'h52dc3dae;
    ram_cell[    2616] = 32'h0;  // 32'h54fa67d7;
    ram_cell[    2617] = 32'h0;  // 32'he93d3ac3;
    ram_cell[    2618] = 32'h0;  // 32'h17d7c09d;
    ram_cell[    2619] = 32'h0;  // 32'h0a220460;
    ram_cell[    2620] = 32'h0;  // 32'h7c9b5f76;
    ram_cell[    2621] = 32'h0;  // 32'h62826d9f;
    ram_cell[    2622] = 32'h0;  // 32'h4a7595fe;
    ram_cell[    2623] = 32'h0;  // 32'h6becb1bd;
    ram_cell[    2624] = 32'h0;  // 32'ha299f633;
    ram_cell[    2625] = 32'h0;  // 32'hfc612425;
    ram_cell[    2626] = 32'h0;  // 32'h994c4c35;
    ram_cell[    2627] = 32'h0;  // 32'hd8ab6e4c;
    ram_cell[    2628] = 32'h0;  // 32'h77ea8e1f;
    ram_cell[    2629] = 32'h0;  // 32'h592a30f9;
    ram_cell[    2630] = 32'h0;  // 32'h1a86ca51;
    ram_cell[    2631] = 32'h0;  // 32'hd9ed115e;
    ram_cell[    2632] = 32'h0;  // 32'hc43fa03d;
    ram_cell[    2633] = 32'h0;  // 32'h1ecbb426;
    ram_cell[    2634] = 32'h0;  // 32'hae1d825e;
    ram_cell[    2635] = 32'h0;  // 32'he8e8e94a;
    ram_cell[    2636] = 32'h0;  // 32'hcd1ed37f;
    ram_cell[    2637] = 32'h0;  // 32'h109bedec;
    ram_cell[    2638] = 32'h0;  // 32'ha573073b;
    ram_cell[    2639] = 32'h0;  // 32'hff54d2b2;
    ram_cell[    2640] = 32'h0;  // 32'h8f6585d1;
    ram_cell[    2641] = 32'h0;  // 32'h85ae83be;
    ram_cell[    2642] = 32'h0;  // 32'h6ace82cd;
    ram_cell[    2643] = 32'h0;  // 32'hd50b00f0;
    ram_cell[    2644] = 32'h0;  // 32'h2a870e93;
    ram_cell[    2645] = 32'h0;  // 32'ha9589bf4;
    ram_cell[    2646] = 32'h0;  // 32'hf29491a5;
    ram_cell[    2647] = 32'h0;  // 32'h28216bbf;
    ram_cell[    2648] = 32'h0;  // 32'h7cdc04c9;
    ram_cell[    2649] = 32'h0;  // 32'hc2e86022;
    ram_cell[    2650] = 32'h0;  // 32'h8e9a0df5;
    ram_cell[    2651] = 32'h0;  // 32'h9221ac39;
    ram_cell[    2652] = 32'h0;  // 32'h3e076ee5;
    ram_cell[    2653] = 32'h0;  // 32'h8f2bd217;
    ram_cell[    2654] = 32'h0;  // 32'h33b0f476;
    ram_cell[    2655] = 32'h0;  // 32'h5de2eb56;
    ram_cell[    2656] = 32'h0;  // 32'h1793425e;
    ram_cell[    2657] = 32'h0;  // 32'h088ef248;
    ram_cell[    2658] = 32'h0;  // 32'h9ff350f1;
    ram_cell[    2659] = 32'h0;  // 32'h9f904b5b;
    ram_cell[    2660] = 32'h0;  // 32'h2ba85e98;
    ram_cell[    2661] = 32'h0;  // 32'h3c76b44f;
    ram_cell[    2662] = 32'h0;  // 32'h6574a77c;
    ram_cell[    2663] = 32'h0;  // 32'h1dd4ef81;
    ram_cell[    2664] = 32'h0;  // 32'h20df96bf;
    ram_cell[    2665] = 32'h0;  // 32'h3b2c2d6f;
    ram_cell[    2666] = 32'h0;  // 32'hecd17ae9;
    ram_cell[    2667] = 32'h0;  // 32'h6ca7bb4d;
    ram_cell[    2668] = 32'h0;  // 32'h8290883e;
    ram_cell[    2669] = 32'h0;  // 32'h3b4873e6;
    ram_cell[    2670] = 32'h0;  // 32'h37ac29ab;
    ram_cell[    2671] = 32'h0;  // 32'h635e6174;
    ram_cell[    2672] = 32'h0;  // 32'h53af2ef1;
    ram_cell[    2673] = 32'h0;  // 32'hba89d551;
    ram_cell[    2674] = 32'h0;  // 32'hb8cfddbd;
    ram_cell[    2675] = 32'h0;  // 32'h8c0b90b1;
    ram_cell[    2676] = 32'h0;  // 32'h6fbb3adf;
    ram_cell[    2677] = 32'h0;  // 32'h7670aa8f;
    ram_cell[    2678] = 32'h0;  // 32'hc16dacbe;
    ram_cell[    2679] = 32'h0;  // 32'h2ee7c6f9;
    ram_cell[    2680] = 32'h0;  // 32'hdb72b33a;
    ram_cell[    2681] = 32'h0;  // 32'h7f71f810;
    ram_cell[    2682] = 32'h0;  // 32'h127e383a;
    ram_cell[    2683] = 32'h0;  // 32'h906ccfab;
    ram_cell[    2684] = 32'h0;  // 32'h8ebbeb7a;
    ram_cell[    2685] = 32'h0;  // 32'h5b163c05;
    ram_cell[    2686] = 32'h0;  // 32'h250cbd92;
    ram_cell[    2687] = 32'h0;  // 32'h5c63e697;
    ram_cell[    2688] = 32'h0;  // 32'hee26471e;
    ram_cell[    2689] = 32'h0;  // 32'h85408c1c;
    ram_cell[    2690] = 32'h0;  // 32'hec984fbe;
    ram_cell[    2691] = 32'h0;  // 32'hde8b37f4;
    ram_cell[    2692] = 32'h0;  // 32'h315f41e0;
    ram_cell[    2693] = 32'h0;  // 32'hf4d6acdb;
    ram_cell[    2694] = 32'h0;  // 32'h616e2d69;
    ram_cell[    2695] = 32'h0;  // 32'h0afb4940;
    ram_cell[    2696] = 32'h0;  // 32'h264b5989;
    ram_cell[    2697] = 32'h0;  // 32'h2a873d24;
    ram_cell[    2698] = 32'h0;  // 32'h732b07e9;
    ram_cell[    2699] = 32'h0;  // 32'h72dc693e;
    ram_cell[    2700] = 32'h0;  // 32'h336a5a1b;
    ram_cell[    2701] = 32'h0;  // 32'h31e3a0bb;
    ram_cell[    2702] = 32'h0;  // 32'hddc02c7d;
    ram_cell[    2703] = 32'h0;  // 32'h0fbeaffe;
    ram_cell[    2704] = 32'h0;  // 32'hc2249ecf;
    ram_cell[    2705] = 32'h0;  // 32'he0e15914;
    ram_cell[    2706] = 32'h0;  // 32'hebb1020b;
    ram_cell[    2707] = 32'h0;  // 32'hc1770d76;
    ram_cell[    2708] = 32'h0;  // 32'ha54b6de7;
    ram_cell[    2709] = 32'h0;  // 32'hc7b7ab5b;
    ram_cell[    2710] = 32'h0;  // 32'heacf1173;
    ram_cell[    2711] = 32'h0;  // 32'h993c0c00;
    ram_cell[    2712] = 32'h0;  // 32'h0bd01f1a;
    ram_cell[    2713] = 32'h0;  // 32'h1f077564;
    ram_cell[    2714] = 32'h0;  // 32'h570e9e17;
    ram_cell[    2715] = 32'h0;  // 32'hcf3ee6e9;
    ram_cell[    2716] = 32'h0;  // 32'h300b5b4b;
    ram_cell[    2717] = 32'h0;  // 32'hf7b3ea5b;
    ram_cell[    2718] = 32'h0;  // 32'hf9cf47f3;
    ram_cell[    2719] = 32'h0;  // 32'hf2d1aeb6;
    ram_cell[    2720] = 32'h0;  // 32'h8da4b1cf;
    ram_cell[    2721] = 32'h0;  // 32'ha36dc5f5;
    ram_cell[    2722] = 32'h0;  // 32'h25b1d246;
    ram_cell[    2723] = 32'h0;  // 32'h0b4a62a8;
    ram_cell[    2724] = 32'h0;  // 32'h59739687;
    ram_cell[    2725] = 32'h0;  // 32'h2ae8251e;
    ram_cell[    2726] = 32'h0;  // 32'ha87b5f52;
    ram_cell[    2727] = 32'h0;  // 32'hf4c01231;
    ram_cell[    2728] = 32'h0;  // 32'hfda6510c;
    ram_cell[    2729] = 32'h0;  // 32'h76586384;
    ram_cell[    2730] = 32'h0;  // 32'hf855fe12;
    ram_cell[    2731] = 32'h0;  // 32'h0e70e5d7;
    ram_cell[    2732] = 32'h0;  // 32'hbb62f42e;
    ram_cell[    2733] = 32'h0;  // 32'hf1eca068;
    ram_cell[    2734] = 32'h0;  // 32'h44e178a1;
    ram_cell[    2735] = 32'h0;  // 32'hfba4c830;
    ram_cell[    2736] = 32'h0;  // 32'h13674118;
    ram_cell[    2737] = 32'h0;  // 32'h2a9f4c9c;
    ram_cell[    2738] = 32'h0;  // 32'h57aa2145;
    ram_cell[    2739] = 32'h0;  // 32'h34994e2d;
    ram_cell[    2740] = 32'h0;  // 32'h89b308cb;
    ram_cell[    2741] = 32'h0;  // 32'he1c23323;
    ram_cell[    2742] = 32'h0;  // 32'hf538c190;
    ram_cell[    2743] = 32'h0;  // 32'h3712b7c8;
    ram_cell[    2744] = 32'h0;  // 32'hdb5481d1;
    ram_cell[    2745] = 32'h0;  // 32'h45b0a7f9;
    ram_cell[    2746] = 32'h0;  // 32'hf00d22b4;
    ram_cell[    2747] = 32'h0;  // 32'h755bdf47;
    ram_cell[    2748] = 32'h0;  // 32'hd4ec4b82;
    ram_cell[    2749] = 32'h0;  // 32'h5804f036;
    ram_cell[    2750] = 32'h0;  // 32'hce800eaa;
    ram_cell[    2751] = 32'h0;  // 32'hee3b747e;
    ram_cell[    2752] = 32'h0;  // 32'hcbb0421e;
    ram_cell[    2753] = 32'h0;  // 32'hc2c6cf55;
    ram_cell[    2754] = 32'h0;  // 32'h2bbf7c89;
    ram_cell[    2755] = 32'h0;  // 32'ha4b35a8f;
    ram_cell[    2756] = 32'h0;  // 32'hbdbee26f;
    ram_cell[    2757] = 32'h0;  // 32'h2a3051ac;
    ram_cell[    2758] = 32'h0;  // 32'h57268771;
    ram_cell[    2759] = 32'h0;  // 32'he0c3fe76;
    ram_cell[    2760] = 32'h0;  // 32'h07a0ac95;
    ram_cell[    2761] = 32'h0;  // 32'h2c8629f4;
    ram_cell[    2762] = 32'h0;  // 32'had5edee4;
    ram_cell[    2763] = 32'h0;  // 32'h4a2a50df;
    ram_cell[    2764] = 32'h0;  // 32'h8c2685d2;
    ram_cell[    2765] = 32'h0;  // 32'h6a46dd02;
    ram_cell[    2766] = 32'h0;  // 32'h329b22ef;
    ram_cell[    2767] = 32'h0;  // 32'hbcf9c3b6;
    ram_cell[    2768] = 32'h0;  // 32'h3cb5f986;
    ram_cell[    2769] = 32'h0;  // 32'h421d06fa;
    ram_cell[    2770] = 32'h0;  // 32'h792135e8;
    ram_cell[    2771] = 32'h0;  // 32'h38980f66;
    ram_cell[    2772] = 32'h0;  // 32'hd4b2cf1b;
    ram_cell[    2773] = 32'h0;  // 32'h6606b5e2;
    ram_cell[    2774] = 32'h0;  // 32'h24e34cb9;
    ram_cell[    2775] = 32'h0;  // 32'h81144392;
    ram_cell[    2776] = 32'h0;  // 32'h53280b09;
    ram_cell[    2777] = 32'h0;  // 32'h81ec72e2;
    ram_cell[    2778] = 32'h0;  // 32'h7124d61a;
    ram_cell[    2779] = 32'h0;  // 32'he7d93303;
    ram_cell[    2780] = 32'h0;  // 32'hceff288d;
    ram_cell[    2781] = 32'h0;  // 32'h26bdf16e;
    ram_cell[    2782] = 32'h0;  // 32'h0eafab8c;
    ram_cell[    2783] = 32'h0;  // 32'h54c4957e;
    ram_cell[    2784] = 32'h0;  // 32'h5e87a70a;
    ram_cell[    2785] = 32'h0;  // 32'h34a27ee6;
    ram_cell[    2786] = 32'h0;  // 32'ha77784b7;
    ram_cell[    2787] = 32'h0;  // 32'h629d18bc;
    ram_cell[    2788] = 32'h0;  // 32'h8ace2495;
    ram_cell[    2789] = 32'h0;  // 32'h407358cc;
    ram_cell[    2790] = 32'h0;  // 32'hcab61ff6;
    ram_cell[    2791] = 32'h0;  // 32'h426e7024;
    ram_cell[    2792] = 32'h0;  // 32'h57b15b3d;
    ram_cell[    2793] = 32'h0;  // 32'hc3705f94;
    ram_cell[    2794] = 32'h0;  // 32'he55a8489;
    ram_cell[    2795] = 32'h0;  // 32'h970fe328;
    ram_cell[    2796] = 32'h0;  // 32'ha510eb04;
    ram_cell[    2797] = 32'h0;  // 32'h8f20f7e0;
    ram_cell[    2798] = 32'h0;  // 32'h5c6ca072;
    ram_cell[    2799] = 32'h0;  // 32'h0dae7443;
    ram_cell[    2800] = 32'h0;  // 32'h4aafd3de;
    ram_cell[    2801] = 32'h0;  // 32'h1a406189;
    ram_cell[    2802] = 32'h0;  // 32'h7f4778e8;
    ram_cell[    2803] = 32'h0;  // 32'h97a7aa0d;
    ram_cell[    2804] = 32'h0;  // 32'h8f7ee411;
    ram_cell[    2805] = 32'h0;  // 32'hee0d9020;
    ram_cell[    2806] = 32'h0;  // 32'h073a4351;
    ram_cell[    2807] = 32'h0;  // 32'h5d3b29de;
    ram_cell[    2808] = 32'h0;  // 32'hf9cff5c6;
    ram_cell[    2809] = 32'h0;  // 32'h499d3dfe;
    ram_cell[    2810] = 32'h0;  // 32'h1f355c61;
    ram_cell[    2811] = 32'h0;  // 32'hf3018056;
    ram_cell[    2812] = 32'h0;  // 32'hdb1d60ab;
    ram_cell[    2813] = 32'h0;  // 32'h5a97ba5f;
    ram_cell[    2814] = 32'h0;  // 32'h4b6648a7;
    ram_cell[    2815] = 32'h0;  // 32'h3baac616;
    ram_cell[    2816] = 32'h0;  // 32'hb8b13b77;
    ram_cell[    2817] = 32'h0;  // 32'h2f19835b;
    ram_cell[    2818] = 32'h0;  // 32'h8e66b0d4;
    ram_cell[    2819] = 32'h0;  // 32'h5828ec0d;
    ram_cell[    2820] = 32'h0;  // 32'he2ed2596;
    ram_cell[    2821] = 32'h0;  // 32'h2cfbd8de;
    ram_cell[    2822] = 32'h0;  // 32'h41a9ef36;
    ram_cell[    2823] = 32'h0;  // 32'h1fa0f3b1;
    ram_cell[    2824] = 32'h0;  // 32'hf764703c;
    ram_cell[    2825] = 32'h0;  // 32'hd13d66d7;
    ram_cell[    2826] = 32'h0;  // 32'h56898b31;
    ram_cell[    2827] = 32'h0;  // 32'he05721fe;
    ram_cell[    2828] = 32'h0;  // 32'h77b469a8;
    ram_cell[    2829] = 32'h0;  // 32'ha7ef4ef4;
    ram_cell[    2830] = 32'h0;  // 32'hf77d4969;
    ram_cell[    2831] = 32'h0;  // 32'h17f70bbe;
    ram_cell[    2832] = 32'h0;  // 32'hfb02ec49;
    ram_cell[    2833] = 32'h0;  // 32'h55985d89;
    ram_cell[    2834] = 32'h0;  // 32'hca58dbc8;
    ram_cell[    2835] = 32'h0;  // 32'h7eea33d9;
    ram_cell[    2836] = 32'h0;  // 32'h92b112ed;
    ram_cell[    2837] = 32'h0;  // 32'h5a1d4dd3;
    ram_cell[    2838] = 32'h0;  // 32'h36a6d419;
    ram_cell[    2839] = 32'h0;  // 32'h83a78aeb;
    ram_cell[    2840] = 32'h0;  // 32'hbf24de51;
    ram_cell[    2841] = 32'h0;  // 32'h311b3746;
    ram_cell[    2842] = 32'h0;  // 32'h41c56550;
    ram_cell[    2843] = 32'h0;  // 32'h145f617f;
    ram_cell[    2844] = 32'h0;  // 32'h51aa1200;
    ram_cell[    2845] = 32'h0;  // 32'h086c49ed;
    ram_cell[    2846] = 32'h0;  // 32'hd7705bc4;
    ram_cell[    2847] = 32'h0;  // 32'h2b00b30e;
    ram_cell[    2848] = 32'h0;  // 32'h326fe56c;
    ram_cell[    2849] = 32'h0;  // 32'h4c4761c6;
    ram_cell[    2850] = 32'h0;  // 32'hc149bf85;
    ram_cell[    2851] = 32'h0;  // 32'h796a5bfe;
    ram_cell[    2852] = 32'h0;  // 32'hcc89bf48;
    ram_cell[    2853] = 32'h0;  // 32'h99349aa3;
    ram_cell[    2854] = 32'h0;  // 32'hb5a9e349;
    ram_cell[    2855] = 32'h0;  // 32'hca9c96bd;
    ram_cell[    2856] = 32'h0;  // 32'h4182d07e;
    ram_cell[    2857] = 32'h0;  // 32'h84597783;
    ram_cell[    2858] = 32'h0;  // 32'h9a4b684f;
    ram_cell[    2859] = 32'h0;  // 32'hb827da28;
    ram_cell[    2860] = 32'h0;  // 32'hd233cc77;
    ram_cell[    2861] = 32'h0;  // 32'h67d1a8cf;
    ram_cell[    2862] = 32'h0;  // 32'hcc1a22d7;
    ram_cell[    2863] = 32'h0;  // 32'h2ab886f1;
    ram_cell[    2864] = 32'h0;  // 32'h78c75b11;
    ram_cell[    2865] = 32'h0;  // 32'h4e161428;
    ram_cell[    2866] = 32'h0;  // 32'h3d564da6;
    ram_cell[    2867] = 32'h0;  // 32'h4c5e7dd7;
    ram_cell[    2868] = 32'h0;  // 32'hb9e1412e;
    ram_cell[    2869] = 32'h0;  // 32'h45385306;
    ram_cell[    2870] = 32'h0;  // 32'h6ebda369;
    ram_cell[    2871] = 32'h0;  // 32'h277457a6;
    ram_cell[    2872] = 32'h0;  // 32'he5a1cc3d;
    ram_cell[    2873] = 32'h0;  // 32'h9e9409cd;
    ram_cell[    2874] = 32'h0;  // 32'h40a46bf8;
    ram_cell[    2875] = 32'h0;  // 32'hd164958f;
    ram_cell[    2876] = 32'h0;  // 32'ha8b60e33;
    ram_cell[    2877] = 32'h0;  // 32'h82e9c92c;
    ram_cell[    2878] = 32'h0;  // 32'ha5c5ca36;
    ram_cell[    2879] = 32'h0;  // 32'heb1a787f;
    ram_cell[    2880] = 32'h0;  // 32'h72e9a96e;
    ram_cell[    2881] = 32'h0;  // 32'h1b96ea7c;
    ram_cell[    2882] = 32'h0;  // 32'h324e3ee5;
    ram_cell[    2883] = 32'h0;  // 32'hfaa725a0;
    ram_cell[    2884] = 32'h0;  // 32'h3cd02b76;
    ram_cell[    2885] = 32'h0;  // 32'h74ea7cfb;
    ram_cell[    2886] = 32'h0;  // 32'h3f6e6924;
    ram_cell[    2887] = 32'h0;  // 32'hdf765b4d;
    ram_cell[    2888] = 32'h0;  // 32'hdc2120f6;
    ram_cell[    2889] = 32'h0;  // 32'h4c7b0150;
    ram_cell[    2890] = 32'h0;  // 32'h5f5d83a4;
    ram_cell[    2891] = 32'h0;  // 32'h1e6f79b7;
    ram_cell[    2892] = 32'h0;  // 32'h82f41010;
    ram_cell[    2893] = 32'h0;  // 32'h0164c986;
    ram_cell[    2894] = 32'h0;  // 32'h762eb2ad;
    ram_cell[    2895] = 32'h0;  // 32'hb7a870d1;
    ram_cell[    2896] = 32'h0;  // 32'he261e2ed;
    ram_cell[    2897] = 32'h0;  // 32'h46a603ab;
    ram_cell[    2898] = 32'h0;  // 32'h40c6e96c;
    ram_cell[    2899] = 32'h0;  // 32'hda138b64;
    ram_cell[    2900] = 32'h0;  // 32'hdb2c24d6;
    ram_cell[    2901] = 32'h0;  // 32'heef64c8d;
    ram_cell[    2902] = 32'h0;  // 32'h47b97bcb;
    ram_cell[    2903] = 32'h0;  // 32'h41a8f66f;
    ram_cell[    2904] = 32'h0;  // 32'h31c88517;
    ram_cell[    2905] = 32'h0;  // 32'h91211423;
    ram_cell[    2906] = 32'h0;  // 32'h203fb6ed;
    ram_cell[    2907] = 32'h0;  // 32'h5347fd65;
    ram_cell[    2908] = 32'h0;  // 32'h73007466;
    ram_cell[    2909] = 32'h0;  // 32'h147d2324;
    ram_cell[    2910] = 32'h0;  // 32'hc28e1098;
    ram_cell[    2911] = 32'h0;  // 32'ha30ef78a;
    ram_cell[    2912] = 32'h0;  // 32'hd2ae5a5d;
    ram_cell[    2913] = 32'h0;  // 32'h1921f109;
    ram_cell[    2914] = 32'h0;  // 32'h163aeded;
    ram_cell[    2915] = 32'h0;  // 32'h1e539fd5;
    ram_cell[    2916] = 32'h0;  // 32'h89d2800f;
    ram_cell[    2917] = 32'h0;  // 32'h0e3c6855;
    ram_cell[    2918] = 32'h0;  // 32'hb756b5ba;
    ram_cell[    2919] = 32'h0;  // 32'hed7eb7eb;
    ram_cell[    2920] = 32'h0;  // 32'he967c9ff;
    ram_cell[    2921] = 32'h0;  // 32'h4bd2e344;
    ram_cell[    2922] = 32'h0;  // 32'h9ddcb37a;
    ram_cell[    2923] = 32'h0;  // 32'hb5492243;
    ram_cell[    2924] = 32'h0;  // 32'h13415585;
    ram_cell[    2925] = 32'h0;  // 32'h7f801540;
    ram_cell[    2926] = 32'h0;  // 32'he107ca17;
    ram_cell[    2927] = 32'h0;  // 32'hfedcaede;
    ram_cell[    2928] = 32'h0;  // 32'hdda0e2f8;
    ram_cell[    2929] = 32'h0;  // 32'h78e0ce3d;
    ram_cell[    2930] = 32'h0;  // 32'h6bacd6a0;
    ram_cell[    2931] = 32'h0;  // 32'hc7a38045;
    ram_cell[    2932] = 32'h0;  // 32'h05b63291;
    ram_cell[    2933] = 32'h0;  // 32'h432f5591;
    ram_cell[    2934] = 32'h0;  // 32'h25cad3ce;
    ram_cell[    2935] = 32'h0;  // 32'h0ccbb7c5;
    ram_cell[    2936] = 32'h0;  // 32'hf6d88f3e;
    ram_cell[    2937] = 32'h0;  // 32'h61c9ade7;
    ram_cell[    2938] = 32'h0;  // 32'hc6bf49c5;
    ram_cell[    2939] = 32'h0;  // 32'h9bbd6581;
    ram_cell[    2940] = 32'h0;  // 32'h4e4ed922;
    ram_cell[    2941] = 32'h0;  // 32'hd076f395;
    ram_cell[    2942] = 32'h0;  // 32'h137dc603;
    ram_cell[    2943] = 32'h0;  // 32'h76273bf8;
    ram_cell[    2944] = 32'h0;  // 32'h1636a1fe;
    ram_cell[    2945] = 32'h0;  // 32'h8f8c12d8;
    ram_cell[    2946] = 32'h0;  // 32'hfa6837a7;
    ram_cell[    2947] = 32'h0;  // 32'h011aba09;
    ram_cell[    2948] = 32'h0;  // 32'h64d66d00;
    ram_cell[    2949] = 32'h0;  // 32'h430c049d;
    ram_cell[    2950] = 32'h0;  // 32'hcd1bf29c;
    ram_cell[    2951] = 32'h0;  // 32'h29c280e6;
    ram_cell[    2952] = 32'h0;  // 32'h84f0c0c1;
    ram_cell[    2953] = 32'h0;  // 32'hf3204342;
    ram_cell[    2954] = 32'h0;  // 32'h16cd6aba;
    ram_cell[    2955] = 32'h0;  // 32'h6ebcff0b;
    ram_cell[    2956] = 32'h0;  // 32'h04ad897e;
    ram_cell[    2957] = 32'h0;  // 32'hda3a6d36;
    ram_cell[    2958] = 32'h0;  // 32'hc30a7a9a;
    ram_cell[    2959] = 32'h0;  // 32'h6c2ab6cb;
    ram_cell[    2960] = 32'h0;  // 32'h00b19cd7;
    ram_cell[    2961] = 32'h0;  // 32'h95d3d73e;
    ram_cell[    2962] = 32'h0;  // 32'h680a61b8;
    ram_cell[    2963] = 32'h0;  // 32'h5bfd23f1;
    ram_cell[    2964] = 32'h0;  // 32'h1cb53945;
    ram_cell[    2965] = 32'h0;  // 32'h7d1530f5;
    ram_cell[    2966] = 32'h0;  // 32'ha81f62b0;
    ram_cell[    2967] = 32'h0;  // 32'h41a4e045;
    ram_cell[    2968] = 32'h0;  // 32'h1043ff35;
    ram_cell[    2969] = 32'h0;  // 32'h249cfd9a;
    ram_cell[    2970] = 32'h0;  // 32'h5df995d1;
    ram_cell[    2971] = 32'h0;  // 32'h7c676803;
    ram_cell[    2972] = 32'h0;  // 32'h196003ac;
    ram_cell[    2973] = 32'h0;  // 32'h07b7ca85;
    ram_cell[    2974] = 32'h0;  // 32'h2cefb2cc;
    ram_cell[    2975] = 32'h0;  // 32'h866f9b46;
    ram_cell[    2976] = 32'h0;  // 32'h99cefbd8;
    ram_cell[    2977] = 32'h0;  // 32'ha87e683f;
    ram_cell[    2978] = 32'h0;  // 32'h4572c8c5;
    ram_cell[    2979] = 32'h0;  // 32'haa99c34b;
    ram_cell[    2980] = 32'h0;  // 32'hba82ee53;
    ram_cell[    2981] = 32'h0;  // 32'h786e0ce4;
    ram_cell[    2982] = 32'h0;  // 32'ha9f036df;
    ram_cell[    2983] = 32'h0;  // 32'h730673c7;
    ram_cell[    2984] = 32'h0;  // 32'hc6e560c3;
    ram_cell[    2985] = 32'h0;  // 32'hde63ce91;
    ram_cell[    2986] = 32'h0;  // 32'h4a8cfffe;
    ram_cell[    2987] = 32'h0;  // 32'h04cc3e4e;
    ram_cell[    2988] = 32'h0;  // 32'hb7083eec;
    ram_cell[    2989] = 32'h0;  // 32'h0e154ffd;
    ram_cell[    2990] = 32'h0;  // 32'h5292e04f;
    ram_cell[    2991] = 32'h0;  // 32'h1d34e080;
    ram_cell[    2992] = 32'h0;  // 32'ha8d50e4a;
    ram_cell[    2993] = 32'h0;  // 32'h67ad4aa0;
    ram_cell[    2994] = 32'h0;  // 32'h2076144b;
    ram_cell[    2995] = 32'h0;  // 32'h65bddf1f;
    ram_cell[    2996] = 32'h0;  // 32'hcfa46154;
    ram_cell[    2997] = 32'h0;  // 32'h555e9df0;
    ram_cell[    2998] = 32'h0;  // 32'hfca6141c;
    ram_cell[    2999] = 32'h0;  // 32'h492b7430;
    ram_cell[    3000] = 32'h0;  // 32'h30c925c6;
    ram_cell[    3001] = 32'h0;  // 32'hd0657946;
    ram_cell[    3002] = 32'h0;  // 32'h78534452;
    ram_cell[    3003] = 32'h0;  // 32'h6fd6ad39;
    ram_cell[    3004] = 32'h0;  // 32'h7aba8ee7;
    ram_cell[    3005] = 32'h0;  // 32'hab148a4f;
    ram_cell[    3006] = 32'h0;  // 32'ha31ca83a;
    ram_cell[    3007] = 32'h0;  // 32'hbd9aa46b;
    ram_cell[    3008] = 32'h0;  // 32'h8c83bd40;
    ram_cell[    3009] = 32'h0;  // 32'h9de4eefd;
    ram_cell[    3010] = 32'h0;  // 32'h0d97ef86;
    ram_cell[    3011] = 32'h0;  // 32'h3e2939f2;
    ram_cell[    3012] = 32'h0;  // 32'haaeb994f;
    ram_cell[    3013] = 32'h0;  // 32'hb9a8b0ce;
    ram_cell[    3014] = 32'h0;  // 32'h47fc37c5;
    ram_cell[    3015] = 32'h0;  // 32'hc1cfc18a;
    ram_cell[    3016] = 32'h0;  // 32'he77ba9b2;
    ram_cell[    3017] = 32'h0;  // 32'hb517afce;
    ram_cell[    3018] = 32'h0;  // 32'h029fa9a9;
    ram_cell[    3019] = 32'h0;  // 32'h71f71ef1;
    ram_cell[    3020] = 32'h0;  // 32'h2f421614;
    ram_cell[    3021] = 32'h0;  // 32'h57b1c1da;
    ram_cell[    3022] = 32'h0;  // 32'h49ad5365;
    ram_cell[    3023] = 32'h0;  // 32'h8e348a81;
    ram_cell[    3024] = 32'h0;  // 32'h9152575e;
    ram_cell[    3025] = 32'h0;  // 32'h1783a168;
    ram_cell[    3026] = 32'h0;  // 32'hae9114b9;
    ram_cell[    3027] = 32'h0;  // 32'h700587eb;
    ram_cell[    3028] = 32'h0;  // 32'hca13e7e0;
    ram_cell[    3029] = 32'h0;  // 32'hdee114fa;
    ram_cell[    3030] = 32'h0;  // 32'h23945f69;
    ram_cell[    3031] = 32'h0;  // 32'h122c1a08;
    ram_cell[    3032] = 32'h0;  // 32'hcc3480a1;
    ram_cell[    3033] = 32'h0;  // 32'hf206c04b;
    ram_cell[    3034] = 32'h0;  // 32'h2b784d1d;
    ram_cell[    3035] = 32'h0;  // 32'h7a6d84c8;
    ram_cell[    3036] = 32'h0;  // 32'h76a12bfa;
    ram_cell[    3037] = 32'h0;  // 32'hdce03c57;
    ram_cell[    3038] = 32'h0;  // 32'h3e9632cd;
    ram_cell[    3039] = 32'h0;  // 32'h494f9b7b;
    ram_cell[    3040] = 32'h0;  // 32'hb02a0dab;
    ram_cell[    3041] = 32'h0;  // 32'hd723b364;
    ram_cell[    3042] = 32'h0;  // 32'h41af993c;
    ram_cell[    3043] = 32'h0;  // 32'h67916bea;
    ram_cell[    3044] = 32'h0;  // 32'h3957a74a;
    ram_cell[    3045] = 32'h0;  // 32'hc5e8d33f;
    ram_cell[    3046] = 32'h0;  // 32'h190d6b01;
    ram_cell[    3047] = 32'h0;  // 32'hf469c4d8;
    ram_cell[    3048] = 32'h0;  // 32'ha6d5ba81;
    ram_cell[    3049] = 32'h0;  // 32'h16d0d02e;
    ram_cell[    3050] = 32'h0;  // 32'hc15c41e2;
    ram_cell[    3051] = 32'h0;  // 32'h6ea3bbcd;
    ram_cell[    3052] = 32'h0;  // 32'hf4a67044;
    ram_cell[    3053] = 32'h0;  // 32'he816289e;
    ram_cell[    3054] = 32'h0;  // 32'h23163e3f;
    ram_cell[    3055] = 32'h0;  // 32'h28e40ea1;
    ram_cell[    3056] = 32'h0;  // 32'h7df23376;
    ram_cell[    3057] = 32'h0;  // 32'hff971512;
    ram_cell[    3058] = 32'h0;  // 32'h7a48fb49;
    ram_cell[    3059] = 32'h0;  // 32'h82723c8e;
    ram_cell[    3060] = 32'h0;  // 32'h0a8bf980;
    ram_cell[    3061] = 32'h0;  // 32'h2171e7bc;
    ram_cell[    3062] = 32'h0;  // 32'h1c8acb8a;
    ram_cell[    3063] = 32'h0;  // 32'h7eba523a;
    ram_cell[    3064] = 32'h0;  // 32'hac2f3804;
    ram_cell[    3065] = 32'h0;  // 32'h843ec8e2;
    ram_cell[    3066] = 32'h0;  // 32'hbaa03218;
    ram_cell[    3067] = 32'h0;  // 32'hef15dd3e;
    ram_cell[    3068] = 32'h0;  // 32'hd72a2677;
    ram_cell[    3069] = 32'h0;  // 32'h4e849731;
    ram_cell[    3070] = 32'h0;  // 32'hb67ac32a;
    ram_cell[    3071] = 32'h0;  // 32'h8b6ff80d;
    ram_cell[    3072] = 32'h0;  // 32'h4febc3c7;
    ram_cell[    3073] = 32'h0;  // 32'hd259edc5;
    ram_cell[    3074] = 32'h0;  // 32'hc3383e4b;
    ram_cell[    3075] = 32'h0;  // 32'h7daecb89;
    ram_cell[    3076] = 32'h0;  // 32'h5649541e;
    ram_cell[    3077] = 32'h0;  // 32'hca281bee;
    ram_cell[    3078] = 32'h0;  // 32'h5fd6836a;
    ram_cell[    3079] = 32'h0;  // 32'h6075ada6;
    ram_cell[    3080] = 32'h0;  // 32'h14b362fb;
    ram_cell[    3081] = 32'h0;  // 32'hac43908f;
    ram_cell[    3082] = 32'h0;  // 32'hf01beb5d;
    ram_cell[    3083] = 32'h0;  // 32'hfe120fc0;
    ram_cell[    3084] = 32'h0;  // 32'h47a2d1b7;
    ram_cell[    3085] = 32'h0;  // 32'h74fbfb9b;
    ram_cell[    3086] = 32'h0;  // 32'hb79a8cb8;
    ram_cell[    3087] = 32'h0;  // 32'h66f66495;
    ram_cell[    3088] = 32'h0;  // 32'hf8ce8f28;
    ram_cell[    3089] = 32'h0;  // 32'h871dc7f5;
    ram_cell[    3090] = 32'h0;  // 32'hcc0e6022;
    ram_cell[    3091] = 32'h0;  // 32'h5ba0416c;
    ram_cell[    3092] = 32'h0;  // 32'h5931f6b5;
    ram_cell[    3093] = 32'h0;  // 32'h033eea6c;
    ram_cell[    3094] = 32'h0;  // 32'h89446c5e;
    ram_cell[    3095] = 32'h0;  // 32'hd7e530e2;
    ram_cell[    3096] = 32'h0;  // 32'h8ba113bd;
    ram_cell[    3097] = 32'h0;  // 32'h4b897f4c;
    ram_cell[    3098] = 32'h0;  // 32'he013d11f;
    ram_cell[    3099] = 32'h0;  // 32'hf046f67a;
    ram_cell[    3100] = 32'h0;  // 32'h7d74279c;
    ram_cell[    3101] = 32'h0;  // 32'he7e2df16;
    ram_cell[    3102] = 32'h0;  // 32'h4d51aaab;
    ram_cell[    3103] = 32'h0;  // 32'h68a9bfcf;
    ram_cell[    3104] = 32'h0;  // 32'hb18b9a4d;
    ram_cell[    3105] = 32'h0;  // 32'h829c435e;
    ram_cell[    3106] = 32'h0;  // 32'hd5886206;
    ram_cell[    3107] = 32'h0;  // 32'h5ccea4d9;
    ram_cell[    3108] = 32'h0;  // 32'h5694b4f6;
    ram_cell[    3109] = 32'h0;  // 32'ha391ebce;
    ram_cell[    3110] = 32'h0;  // 32'ha226c189;
    ram_cell[    3111] = 32'h0;  // 32'h2d5f19de;
    ram_cell[    3112] = 32'h0;  // 32'h16254bf8;
    ram_cell[    3113] = 32'h0;  // 32'h47173f16;
    ram_cell[    3114] = 32'h0;  // 32'habe55606;
    ram_cell[    3115] = 32'h0;  // 32'h1df7687f;
    ram_cell[    3116] = 32'h0;  // 32'hc48dd282;
    ram_cell[    3117] = 32'h0;  // 32'hf2689b97;
    ram_cell[    3118] = 32'h0;  // 32'h3db1df8b;
    ram_cell[    3119] = 32'h0;  // 32'hdc80706b;
    ram_cell[    3120] = 32'h0;  // 32'hfa7e7d1f;
    ram_cell[    3121] = 32'h0;  // 32'hb98ed67a;
    ram_cell[    3122] = 32'h0;  // 32'h5442f60c;
    ram_cell[    3123] = 32'h0;  // 32'hf3ed44ef;
    ram_cell[    3124] = 32'h0;  // 32'h42097f3c;
    ram_cell[    3125] = 32'h0;  // 32'h5d0837a3;
    ram_cell[    3126] = 32'h0;  // 32'h482c38d3;
    ram_cell[    3127] = 32'h0;  // 32'h05b1caf7;
    ram_cell[    3128] = 32'h0;  // 32'hb3e86edc;
    ram_cell[    3129] = 32'h0;  // 32'h900eb9c5;
    ram_cell[    3130] = 32'h0;  // 32'h6ba3b5c5;
    ram_cell[    3131] = 32'h0;  // 32'h98976d49;
    ram_cell[    3132] = 32'h0;  // 32'haed028ce;
    ram_cell[    3133] = 32'h0;  // 32'hd70fa7c3;
    ram_cell[    3134] = 32'h0;  // 32'h95b47275;
    ram_cell[    3135] = 32'h0;  // 32'h1e3b52aa;
    ram_cell[    3136] = 32'h0;  // 32'h79234fbc;
    ram_cell[    3137] = 32'h0;  // 32'h95ebad84;
    ram_cell[    3138] = 32'h0;  // 32'h915e5472;
    ram_cell[    3139] = 32'h0;  // 32'h02ac820d;
    ram_cell[    3140] = 32'h0;  // 32'h19a11d7e;
    ram_cell[    3141] = 32'h0;  // 32'h197133bf;
    ram_cell[    3142] = 32'h0;  // 32'h667c054f;
    ram_cell[    3143] = 32'h0;  // 32'hfd9c9d18;
    ram_cell[    3144] = 32'h0;  // 32'h3f4efc04;
    ram_cell[    3145] = 32'h0;  // 32'hc2c20149;
    ram_cell[    3146] = 32'h0;  // 32'hbaa0bc2f;
    ram_cell[    3147] = 32'h0;  // 32'h41c442a0;
    ram_cell[    3148] = 32'h0;  // 32'h7f84eaab;
    ram_cell[    3149] = 32'h0;  // 32'hdcdcd0a9;
    ram_cell[    3150] = 32'h0;  // 32'h860ca423;
    ram_cell[    3151] = 32'h0;  // 32'hf013d67a;
    ram_cell[    3152] = 32'h0;  // 32'h6a6a5c31;
    ram_cell[    3153] = 32'h0;  // 32'hd8744995;
    ram_cell[    3154] = 32'h0;  // 32'hf8025a79;
    ram_cell[    3155] = 32'h0;  // 32'h03af2876;
    ram_cell[    3156] = 32'h0;  // 32'h9628797d;
    ram_cell[    3157] = 32'h0;  // 32'h09500865;
    ram_cell[    3158] = 32'h0;  // 32'h68780c80;
    ram_cell[    3159] = 32'h0;  // 32'h799b59eb;
    ram_cell[    3160] = 32'h0;  // 32'h0fdc8c9d;
    ram_cell[    3161] = 32'h0;  // 32'h7eae8307;
    ram_cell[    3162] = 32'h0;  // 32'ha55ed484;
    ram_cell[    3163] = 32'h0;  // 32'h5ed5693c;
    ram_cell[    3164] = 32'h0;  // 32'h43e808f7;
    ram_cell[    3165] = 32'h0;  // 32'h6d6c76ec;
    ram_cell[    3166] = 32'h0;  // 32'hf0052b5b;
    ram_cell[    3167] = 32'h0;  // 32'hc088e095;
    ram_cell[    3168] = 32'h0;  // 32'hf329cbf7;
    ram_cell[    3169] = 32'h0;  // 32'he323bdd8;
    ram_cell[    3170] = 32'h0;  // 32'h016f49f4;
    ram_cell[    3171] = 32'h0;  // 32'h94290d2d;
    ram_cell[    3172] = 32'h0;  // 32'h4a122194;
    ram_cell[    3173] = 32'h0;  // 32'hc51b0aa8;
    ram_cell[    3174] = 32'h0;  // 32'h1b0babb2;
    ram_cell[    3175] = 32'h0;  // 32'h61138a04;
    ram_cell[    3176] = 32'h0;  // 32'hdd7deacc;
    ram_cell[    3177] = 32'h0;  // 32'ha9b36932;
    ram_cell[    3178] = 32'h0;  // 32'h8e44b93d;
    ram_cell[    3179] = 32'h0;  // 32'hd14954fb;
    ram_cell[    3180] = 32'h0;  // 32'hea919b8b;
    ram_cell[    3181] = 32'h0;  // 32'hee042d83;
    ram_cell[    3182] = 32'h0;  // 32'he80a8297;
    ram_cell[    3183] = 32'h0;  // 32'ha614b569;
    ram_cell[    3184] = 32'h0;  // 32'h7d1fa476;
    ram_cell[    3185] = 32'h0;  // 32'hfbe5571b;
    ram_cell[    3186] = 32'h0;  // 32'h16156c85;
    ram_cell[    3187] = 32'h0;  // 32'hab8f2741;
    ram_cell[    3188] = 32'h0;  // 32'h0f111977;
    ram_cell[    3189] = 32'h0;  // 32'h5ce59d4d;
    ram_cell[    3190] = 32'h0;  // 32'hb370d301;
    ram_cell[    3191] = 32'h0;  // 32'h406c752a;
    ram_cell[    3192] = 32'h0;  // 32'hdba22599;
    ram_cell[    3193] = 32'h0;  // 32'hd5ff5f0f;
    ram_cell[    3194] = 32'h0;  // 32'h50c4595b;
    ram_cell[    3195] = 32'h0;  // 32'hd7dc2f92;
    ram_cell[    3196] = 32'h0;  // 32'hcdd519c9;
    ram_cell[    3197] = 32'h0;  // 32'h3453c3d2;
    ram_cell[    3198] = 32'h0;  // 32'h2035de3a;
    ram_cell[    3199] = 32'h0;  // 32'h581539a4;
    ram_cell[    3200] = 32'h0;  // 32'hd68a6345;
    ram_cell[    3201] = 32'h0;  // 32'h456bf161;
    ram_cell[    3202] = 32'h0;  // 32'h536ea92e;
    ram_cell[    3203] = 32'h0;  // 32'he497d487;
    ram_cell[    3204] = 32'h0;  // 32'hf2fb7da3;
    ram_cell[    3205] = 32'h0;  // 32'he84142ad;
    ram_cell[    3206] = 32'h0;  // 32'h9d624b2f;
    ram_cell[    3207] = 32'h0;  // 32'h8c5817d9;
    ram_cell[    3208] = 32'h0;  // 32'hcf205ca1;
    ram_cell[    3209] = 32'h0;  // 32'hf4d23537;
    ram_cell[    3210] = 32'h0;  // 32'hcf7aad54;
    ram_cell[    3211] = 32'h0;  // 32'hec6aca4c;
    ram_cell[    3212] = 32'h0;  // 32'hd00be10c;
    ram_cell[    3213] = 32'h0;  // 32'hf2f64fd4;
    ram_cell[    3214] = 32'h0;  // 32'hd19c9098;
    ram_cell[    3215] = 32'h0;  // 32'hd9a5f6d4;
    ram_cell[    3216] = 32'h0;  // 32'haaebb86f;
    ram_cell[    3217] = 32'h0;  // 32'h29e7c7f0;
    ram_cell[    3218] = 32'h0;  // 32'h426d68d3;
    ram_cell[    3219] = 32'h0;  // 32'hb868cc91;
    ram_cell[    3220] = 32'h0;  // 32'h2522f98d;
    ram_cell[    3221] = 32'h0;  // 32'hc57a4381;
    ram_cell[    3222] = 32'h0;  // 32'h3f92d009;
    ram_cell[    3223] = 32'h0;  // 32'hc9b1cc1d;
    ram_cell[    3224] = 32'h0;  // 32'h3e3b0046;
    ram_cell[    3225] = 32'h0;  // 32'h70593f7e;
    ram_cell[    3226] = 32'h0;  // 32'h28b0d353;
    ram_cell[    3227] = 32'h0;  // 32'h9f39d5b8;
    ram_cell[    3228] = 32'h0;  // 32'h5c3d7dd5;
    ram_cell[    3229] = 32'h0;  // 32'h35950fb3;
    ram_cell[    3230] = 32'h0;  // 32'h2c93a62c;
    ram_cell[    3231] = 32'h0;  // 32'h39526661;
    ram_cell[    3232] = 32'h0;  // 32'h9ccde1cb;
    ram_cell[    3233] = 32'h0;  // 32'he70046a8;
    ram_cell[    3234] = 32'h0;  // 32'h9bf4e60e;
    ram_cell[    3235] = 32'h0;  // 32'h9b6900c5;
    ram_cell[    3236] = 32'h0;  // 32'he749706f;
    ram_cell[    3237] = 32'h0;  // 32'he2aa514c;
    ram_cell[    3238] = 32'h0;  // 32'h544d756e;
    ram_cell[    3239] = 32'h0;  // 32'h1caca216;
    ram_cell[    3240] = 32'h0;  // 32'h431afbb1;
    ram_cell[    3241] = 32'h0;  // 32'h1ed6a012;
    ram_cell[    3242] = 32'h0;  // 32'hec689172;
    ram_cell[    3243] = 32'h0;  // 32'h543ef44b;
    ram_cell[    3244] = 32'h0;  // 32'h110c2c0e;
    ram_cell[    3245] = 32'h0;  // 32'h589f1193;
    ram_cell[    3246] = 32'h0;  // 32'hcc8204d5;
    ram_cell[    3247] = 32'h0;  // 32'h13bf87d1;
    ram_cell[    3248] = 32'h0;  // 32'hdceff8ca;
    ram_cell[    3249] = 32'h0;  // 32'hca9d649b;
    ram_cell[    3250] = 32'h0;  // 32'h7e014b41;
    ram_cell[    3251] = 32'h0;  // 32'hf7ac3dc8;
    ram_cell[    3252] = 32'h0;  // 32'he214c7b1;
    ram_cell[    3253] = 32'h0;  // 32'h37c19d86;
    ram_cell[    3254] = 32'h0;  // 32'h1e4fd24d;
    ram_cell[    3255] = 32'h0;  // 32'ha601362a;
    ram_cell[    3256] = 32'h0;  // 32'hc41b14d3;
    ram_cell[    3257] = 32'h0;  // 32'hcfbc6a17;
    ram_cell[    3258] = 32'h0;  // 32'hb8bd3853;
    ram_cell[    3259] = 32'h0;  // 32'hc0e69aa3;
    ram_cell[    3260] = 32'h0;  // 32'h5e50e87a;
    ram_cell[    3261] = 32'h0;  // 32'h15a46e39;
    ram_cell[    3262] = 32'h0;  // 32'h38feb786;
    ram_cell[    3263] = 32'h0;  // 32'hf26af5a8;
    ram_cell[    3264] = 32'h0;  // 32'hfe52e2b7;
    ram_cell[    3265] = 32'h0;  // 32'h3900da0d;
    ram_cell[    3266] = 32'h0;  // 32'h5d83fb75;
    ram_cell[    3267] = 32'h0;  // 32'he4d14a76;
    ram_cell[    3268] = 32'h0;  // 32'h820eb5de;
    ram_cell[    3269] = 32'h0;  // 32'h86db13a0;
    ram_cell[    3270] = 32'h0;  // 32'h1e7f2c17;
    ram_cell[    3271] = 32'h0;  // 32'h3eab23ba;
    ram_cell[    3272] = 32'h0;  // 32'h13960f37;
    ram_cell[    3273] = 32'h0;  // 32'hcfb92065;
    ram_cell[    3274] = 32'h0;  // 32'ha68fb2aa;
    ram_cell[    3275] = 32'h0;  // 32'ha95b93a1;
    ram_cell[    3276] = 32'h0;  // 32'h15066629;
    ram_cell[    3277] = 32'h0;  // 32'hfb343e2a;
    ram_cell[    3278] = 32'h0;  // 32'h4d814e2e;
    ram_cell[    3279] = 32'h0;  // 32'h5f38f5ba;
    ram_cell[    3280] = 32'h0;  // 32'hc0408d00;
    ram_cell[    3281] = 32'h0;  // 32'h37d60ff5;
    ram_cell[    3282] = 32'h0;  // 32'he25cbe67;
    ram_cell[    3283] = 32'h0;  // 32'hf090457f;
    ram_cell[    3284] = 32'h0;  // 32'h08da63e5;
    ram_cell[    3285] = 32'h0;  // 32'h351a5b82;
    ram_cell[    3286] = 32'h0;  // 32'h4c11961f;
    ram_cell[    3287] = 32'h0;  // 32'h96899b1d;
    ram_cell[    3288] = 32'h0;  // 32'hdd3893fb;
    ram_cell[    3289] = 32'h0;  // 32'h6fd1c47e;
    ram_cell[    3290] = 32'h0;  // 32'h06bb563e;
    ram_cell[    3291] = 32'h0;  // 32'h4ab2f9a3;
    ram_cell[    3292] = 32'h0;  // 32'he6cec71e;
    ram_cell[    3293] = 32'h0;  // 32'hf76b4ded;
    ram_cell[    3294] = 32'h0;  // 32'hb4e92bf6;
    ram_cell[    3295] = 32'h0;  // 32'h05cd748c;
    ram_cell[    3296] = 32'h0;  // 32'hdbf97c84;
    ram_cell[    3297] = 32'h0;  // 32'h4c196449;
    ram_cell[    3298] = 32'h0;  // 32'h4f6d633c;
    ram_cell[    3299] = 32'h0;  // 32'hff5690b1;
    ram_cell[    3300] = 32'h0;  // 32'hf46a8f38;
    ram_cell[    3301] = 32'h0;  // 32'hcba0f0d0;
    ram_cell[    3302] = 32'h0;  // 32'h02ef1e5f;
    ram_cell[    3303] = 32'h0;  // 32'h9bca6d98;
    ram_cell[    3304] = 32'h0;  // 32'h52f39a27;
    ram_cell[    3305] = 32'h0;  // 32'h426679f6;
    ram_cell[    3306] = 32'h0;  // 32'h1b2582ae;
    ram_cell[    3307] = 32'h0;  // 32'hc93a4b55;
    ram_cell[    3308] = 32'h0;  // 32'h6b0dc6e4;
    ram_cell[    3309] = 32'h0;  // 32'h471a1346;
    ram_cell[    3310] = 32'h0;  // 32'h6cd23d7e;
    ram_cell[    3311] = 32'h0;  // 32'h6e4c82dc;
    ram_cell[    3312] = 32'h0;  // 32'h89c557c5;
    ram_cell[    3313] = 32'h0;  // 32'h6b469e6d;
    ram_cell[    3314] = 32'h0;  // 32'h7c16b7e4;
    ram_cell[    3315] = 32'h0;  // 32'hd2351536;
    ram_cell[    3316] = 32'h0;  // 32'h5bdbf0b6;
    ram_cell[    3317] = 32'h0;  // 32'h9a3d8503;
    ram_cell[    3318] = 32'h0;  // 32'h72c7d62f;
    ram_cell[    3319] = 32'h0;  // 32'ha58c8870;
    ram_cell[    3320] = 32'h0;  // 32'ha77e34dc;
    ram_cell[    3321] = 32'h0;  // 32'h112ee9e0;
    ram_cell[    3322] = 32'h0;  // 32'h0f8ede43;
    ram_cell[    3323] = 32'h0;  // 32'h42bc3c6b;
    ram_cell[    3324] = 32'h0;  // 32'h1934bc34;
    ram_cell[    3325] = 32'h0;  // 32'h866b2dca;
    ram_cell[    3326] = 32'h0;  // 32'he29d3c5d;
    ram_cell[    3327] = 32'h0;  // 32'h427f0393;
    ram_cell[    3328] = 32'h0;  // 32'hf5d77f7f;
    ram_cell[    3329] = 32'h0;  // 32'h53a593f9;
    ram_cell[    3330] = 32'h0;  // 32'h6f06fb8f;
    ram_cell[    3331] = 32'h0;  // 32'h41cd7a7c;
    ram_cell[    3332] = 32'h0;  // 32'hb81cfc28;
    ram_cell[    3333] = 32'h0;  // 32'h9be165f3;
    ram_cell[    3334] = 32'h0;  // 32'h9dc7daa5;
    ram_cell[    3335] = 32'h0;  // 32'hb4a97b8e;
    ram_cell[    3336] = 32'h0;  // 32'hc51dd8cd;
    ram_cell[    3337] = 32'h0;  // 32'h9d196be6;
    ram_cell[    3338] = 32'h0;  // 32'h0a8e384f;
    ram_cell[    3339] = 32'h0;  // 32'h53bd9025;
    ram_cell[    3340] = 32'h0;  // 32'he7fbf953;
    ram_cell[    3341] = 32'h0;  // 32'h8a3de30f;
    ram_cell[    3342] = 32'h0;  // 32'h36d2ee91;
    ram_cell[    3343] = 32'h0;  // 32'h4db64b33;
    ram_cell[    3344] = 32'h0;  // 32'h785d1d25;
    ram_cell[    3345] = 32'h0;  // 32'heed94177;
    ram_cell[    3346] = 32'h0;  // 32'h3d2e943a;
    ram_cell[    3347] = 32'h0;  // 32'hfd696855;
    ram_cell[    3348] = 32'h0;  // 32'h3a41d034;
    ram_cell[    3349] = 32'h0;  // 32'h3164bbe1;
    ram_cell[    3350] = 32'h0;  // 32'h63d6598e;
    ram_cell[    3351] = 32'h0;  // 32'h45baac46;
    ram_cell[    3352] = 32'h0;  // 32'h127070de;
    ram_cell[    3353] = 32'h0;  // 32'h0bf9afab;
    ram_cell[    3354] = 32'h0;  // 32'h67ae0d16;
    ram_cell[    3355] = 32'h0;  // 32'h7cd81d3a;
    ram_cell[    3356] = 32'h0;  // 32'h076e6f49;
    ram_cell[    3357] = 32'h0;  // 32'h7c7817f3;
    ram_cell[    3358] = 32'h0;  // 32'hb6944e0e;
    ram_cell[    3359] = 32'h0;  // 32'h66782680;
    ram_cell[    3360] = 32'h0;  // 32'h5a35f0b2;
    ram_cell[    3361] = 32'h0;  // 32'he8d417a0;
    ram_cell[    3362] = 32'h0;  // 32'hb70a3610;
    ram_cell[    3363] = 32'h0;  // 32'h11cac11b;
    ram_cell[    3364] = 32'h0;  // 32'hec784d14;
    ram_cell[    3365] = 32'h0;  // 32'had0c3007;
    ram_cell[    3366] = 32'h0;  // 32'h9ea6c16e;
    ram_cell[    3367] = 32'h0;  // 32'hf599070c;
    ram_cell[    3368] = 32'h0;  // 32'hc747bdbc;
    ram_cell[    3369] = 32'h0;  // 32'ha106af87;
    ram_cell[    3370] = 32'h0;  // 32'h76d0f359;
    ram_cell[    3371] = 32'h0;  // 32'ha339ed60;
    ram_cell[    3372] = 32'h0;  // 32'hdec5f99f;
    ram_cell[    3373] = 32'h0;  // 32'h8f97eae2;
    ram_cell[    3374] = 32'h0;  // 32'had06f27b;
    ram_cell[    3375] = 32'h0;  // 32'ha8c95671;
    ram_cell[    3376] = 32'h0;  // 32'h3e06c58a;
    ram_cell[    3377] = 32'h0;  // 32'h89056cd3;
    ram_cell[    3378] = 32'h0;  // 32'h454c7927;
    ram_cell[    3379] = 32'h0;  // 32'h3fd26312;
    ram_cell[    3380] = 32'h0;  // 32'h0c14f201;
    ram_cell[    3381] = 32'h0;  // 32'h575f6f52;
    ram_cell[    3382] = 32'h0;  // 32'he0ca81ed;
    ram_cell[    3383] = 32'h0;  // 32'h8f80e8de;
    ram_cell[    3384] = 32'h0;  // 32'hdd17913c;
    ram_cell[    3385] = 32'h0;  // 32'h543e89b1;
    ram_cell[    3386] = 32'h0;  // 32'hd0420ed9;
    ram_cell[    3387] = 32'h0;  // 32'head11ae2;
    ram_cell[    3388] = 32'h0;  // 32'hca572ba9;
    ram_cell[    3389] = 32'h0;  // 32'h4cb46772;
    ram_cell[    3390] = 32'h0;  // 32'h8fbf6f62;
    ram_cell[    3391] = 32'h0;  // 32'h30fb333a;
    ram_cell[    3392] = 32'h0;  // 32'h5cc749ce;
    ram_cell[    3393] = 32'h0;  // 32'hce0aa3a6;
    ram_cell[    3394] = 32'h0;  // 32'hdc5a6896;
    ram_cell[    3395] = 32'h0;  // 32'h28ce3208;
    ram_cell[    3396] = 32'h0;  // 32'h5ad93464;
    ram_cell[    3397] = 32'h0;  // 32'h1215244e;
    ram_cell[    3398] = 32'h0;  // 32'hf01bf03e;
    ram_cell[    3399] = 32'h0;  // 32'hd975420f;
    ram_cell[    3400] = 32'h0;  // 32'hbbc836ea;
    ram_cell[    3401] = 32'h0;  // 32'hdd3e1927;
    ram_cell[    3402] = 32'h0;  // 32'hc8fc7e52;
    ram_cell[    3403] = 32'h0;  // 32'hae5b2230;
    ram_cell[    3404] = 32'h0;  // 32'had13432a;
    ram_cell[    3405] = 32'h0;  // 32'h408fd100;
    ram_cell[    3406] = 32'h0;  // 32'ha5ffbe8b;
    ram_cell[    3407] = 32'h0;  // 32'hd1ad57a4;
    ram_cell[    3408] = 32'h0;  // 32'hcbe140a9;
    ram_cell[    3409] = 32'h0;  // 32'h9c1b3011;
    ram_cell[    3410] = 32'h0;  // 32'h579e8c2c;
    ram_cell[    3411] = 32'h0;  // 32'he7b9e47b;
    ram_cell[    3412] = 32'h0;  // 32'hb99e7d15;
    ram_cell[    3413] = 32'h0;  // 32'hd5d562c8;
    ram_cell[    3414] = 32'h0;  // 32'h773c0881;
    ram_cell[    3415] = 32'h0;  // 32'h23058d32;
    ram_cell[    3416] = 32'h0;  // 32'he029d8dc;
    ram_cell[    3417] = 32'h0;  // 32'h05869726;
    ram_cell[    3418] = 32'h0;  // 32'hefccb4b0;
    ram_cell[    3419] = 32'h0;  // 32'h215663cb;
    ram_cell[    3420] = 32'h0;  // 32'h06bf31b3;
    ram_cell[    3421] = 32'h0;  // 32'h339e40d9;
    ram_cell[    3422] = 32'h0;  // 32'hcef10bdf;
    ram_cell[    3423] = 32'h0;  // 32'h3b398b8c;
    ram_cell[    3424] = 32'h0;  // 32'h660df06f;
    ram_cell[    3425] = 32'h0;  // 32'ha7e5e97c;
    ram_cell[    3426] = 32'h0;  // 32'h59feab82;
    ram_cell[    3427] = 32'h0;  // 32'hbd53b427;
    ram_cell[    3428] = 32'h0;  // 32'hfec47551;
    ram_cell[    3429] = 32'h0;  // 32'hb3e9af88;
    ram_cell[    3430] = 32'h0;  // 32'hcd5f33f9;
    ram_cell[    3431] = 32'h0;  // 32'h46c09f1c;
    ram_cell[    3432] = 32'h0;  // 32'h5fdad434;
    ram_cell[    3433] = 32'h0;  // 32'h5917dd8b;
    ram_cell[    3434] = 32'h0;  // 32'h3167de22;
    ram_cell[    3435] = 32'h0;  // 32'h81a0732f;
    ram_cell[    3436] = 32'h0;  // 32'h9d79bce2;
    ram_cell[    3437] = 32'h0;  // 32'h4d6dd83b;
    ram_cell[    3438] = 32'h0;  // 32'h6b0114eb;
    ram_cell[    3439] = 32'h0;  // 32'h63f59847;
    ram_cell[    3440] = 32'h0;  // 32'he46e31eb;
    ram_cell[    3441] = 32'h0;  // 32'h9bb5247c;
    ram_cell[    3442] = 32'h0;  // 32'h063f0558;
    ram_cell[    3443] = 32'h0;  // 32'h88558906;
    ram_cell[    3444] = 32'h0;  // 32'h0a946f5d;
    ram_cell[    3445] = 32'h0;  // 32'h918bf8b4;
    ram_cell[    3446] = 32'h0;  // 32'h94bab6a4;
    ram_cell[    3447] = 32'h0;  // 32'hb96a53f2;
    ram_cell[    3448] = 32'h0;  // 32'hbdb7f7d1;
    ram_cell[    3449] = 32'h0;  // 32'hadb0d647;
    ram_cell[    3450] = 32'h0;  // 32'h4234edc3;
    ram_cell[    3451] = 32'h0;  // 32'h6a22577f;
    ram_cell[    3452] = 32'h0;  // 32'h513d38ea;
    ram_cell[    3453] = 32'h0;  // 32'h3ba9374b;
    ram_cell[    3454] = 32'h0;  // 32'h15797755;
    ram_cell[    3455] = 32'h0;  // 32'h92f3b8a9;
    ram_cell[    3456] = 32'h0;  // 32'h02e02fb8;
    ram_cell[    3457] = 32'h0;  // 32'hdc5c82ad;
    ram_cell[    3458] = 32'h0;  // 32'h1021f806;
    ram_cell[    3459] = 32'h0;  // 32'ha0fd25f9;
    ram_cell[    3460] = 32'h0;  // 32'hd2945078;
    ram_cell[    3461] = 32'h0;  // 32'h8d2727e2;
    ram_cell[    3462] = 32'h0;  // 32'h65553e18;
    ram_cell[    3463] = 32'h0;  // 32'h76faccf4;
    ram_cell[    3464] = 32'h0;  // 32'hbb62e159;
    ram_cell[    3465] = 32'h0;  // 32'h9a57ba84;
    ram_cell[    3466] = 32'h0;  // 32'h96860776;
    ram_cell[    3467] = 32'h0;  // 32'h6fce51f5;
    ram_cell[    3468] = 32'h0;  // 32'h9ff0bbe3;
    ram_cell[    3469] = 32'h0;  // 32'h3100add3;
    ram_cell[    3470] = 32'h0;  // 32'h0aa7131a;
    ram_cell[    3471] = 32'h0;  // 32'h099efb22;
    ram_cell[    3472] = 32'h0;  // 32'ha0b8571e;
    ram_cell[    3473] = 32'h0;  // 32'h780e4fbb;
    ram_cell[    3474] = 32'h0;  // 32'h641f47e0;
    ram_cell[    3475] = 32'h0;  // 32'h95f35cf2;
    ram_cell[    3476] = 32'h0;  // 32'h4b51a56b;
    ram_cell[    3477] = 32'h0;  // 32'h2b149043;
    ram_cell[    3478] = 32'h0;  // 32'h383199a2;
    ram_cell[    3479] = 32'h0;  // 32'hdd07d1ac;
    ram_cell[    3480] = 32'h0;  // 32'ha9cd542c;
    ram_cell[    3481] = 32'h0;  // 32'h14f10886;
    ram_cell[    3482] = 32'h0;  // 32'h18d83c34;
    ram_cell[    3483] = 32'h0;  // 32'h33f07d8a;
    ram_cell[    3484] = 32'h0;  // 32'h3fd58ca4;
    ram_cell[    3485] = 32'h0;  // 32'he325e991;
    ram_cell[    3486] = 32'h0;  // 32'hd8d759fb;
    ram_cell[    3487] = 32'h0;  // 32'h3a68c695;
    ram_cell[    3488] = 32'h0;  // 32'h05ea2870;
    ram_cell[    3489] = 32'h0;  // 32'ha54052d3;
    ram_cell[    3490] = 32'h0;  // 32'h1ee38604;
    ram_cell[    3491] = 32'h0;  // 32'h3bce2325;
    ram_cell[    3492] = 32'h0;  // 32'h3cdcea94;
    ram_cell[    3493] = 32'h0;  // 32'hbc64c812;
    ram_cell[    3494] = 32'h0;  // 32'h3265973d;
    ram_cell[    3495] = 32'h0;  // 32'hae929de1;
    ram_cell[    3496] = 32'h0;  // 32'h46c1cac5;
    ram_cell[    3497] = 32'h0;  // 32'hc404848c;
    ram_cell[    3498] = 32'h0;  // 32'h46c3575d;
    ram_cell[    3499] = 32'h0;  // 32'hf51807b7;
    ram_cell[    3500] = 32'h0;  // 32'h6960db48;
    ram_cell[    3501] = 32'h0;  // 32'hcbcc2ebf;
    ram_cell[    3502] = 32'h0;  // 32'h3ccb72b5;
    ram_cell[    3503] = 32'h0;  // 32'hc03a8c6c;
    ram_cell[    3504] = 32'h0;  // 32'hf2432f2d;
    ram_cell[    3505] = 32'h0;  // 32'hc979123e;
    ram_cell[    3506] = 32'h0;  // 32'h4a74f114;
    ram_cell[    3507] = 32'h0;  // 32'h62dd79ac;
    ram_cell[    3508] = 32'h0;  // 32'h18c6f4cc;
    ram_cell[    3509] = 32'h0;  // 32'h760cbfb3;
    ram_cell[    3510] = 32'h0;  // 32'hd0b43dad;
    ram_cell[    3511] = 32'h0;  // 32'h99ea3ff0;
    ram_cell[    3512] = 32'h0;  // 32'h43a56310;
    ram_cell[    3513] = 32'h0;  // 32'hd3e611c2;
    ram_cell[    3514] = 32'h0;  // 32'h72f12143;
    ram_cell[    3515] = 32'h0;  // 32'h44b9eb21;
    ram_cell[    3516] = 32'h0;  // 32'h1c1bf3da;
    ram_cell[    3517] = 32'h0;  // 32'hbae4bd85;
    ram_cell[    3518] = 32'h0;  // 32'hed87c49e;
    ram_cell[    3519] = 32'h0;  // 32'hb70cdaa8;
    ram_cell[    3520] = 32'h0;  // 32'hbd4f484a;
    ram_cell[    3521] = 32'h0;  // 32'hf7cb16d5;
    ram_cell[    3522] = 32'h0;  // 32'ha8a529dd;
    ram_cell[    3523] = 32'h0;  // 32'hec484934;
    ram_cell[    3524] = 32'h0;  // 32'h236a1789;
    ram_cell[    3525] = 32'h0;  // 32'hf2d315fe;
    ram_cell[    3526] = 32'h0;  // 32'h77f27142;
    ram_cell[    3527] = 32'h0;  // 32'h4f6467b3;
    ram_cell[    3528] = 32'h0;  // 32'h42755bf2;
    ram_cell[    3529] = 32'h0;  // 32'h1598a010;
    ram_cell[    3530] = 32'h0;  // 32'hf9b20446;
    ram_cell[    3531] = 32'h0;  // 32'hd818164d;
    ram_cell[    3532] = 32'h0;  // 32'h69b3ed05;
    ram_cell[    3533] = 32'h0;  // 32'hd66a83b1;
    ram_cell[    3534] = 32'h0;  // 32'h16cb36ed;
    ram_cell[    3535] = 32'h0;  // 32'hda7a7fd3;
    ram_cell[    3536] = 32'h0;  // 32'he1bd4a08;
    ram_cell[    3537] = 32'h0;  // 32'h3720f1a8;
    ram_cell[    3538] = 32'h0;  // 32'h9271cabf;
    ram_cell[    3539] = 32'h0;  // 32'hc5186be7;
    ram_cell[    3540] = 32'h0;  // 32'hfdb244b3;
    ram_cell[    3541] = 32'h0;  // 32'h7b9eca39;
    ram_cell[    3542] = 32'h0;  // 32'hbc1b0643;
    ram_cell[    3543] = 32'h0;  // 32'h176f70a5;
    ram_cell[    3544] = 32'h0;  // 32'h9e1043e7;
    ram_cell[    3545] = 32'h0;  // 32'h058eb40e;
    ram_cell[    3546] = 32'h0;  // 32'hc5804460;
    ram_cell[    3547] = 32'h0;  // 32'hcd355935;
    ram_cell[    3548] = 32'h0;  // 32'ha70e03f3;
    ram_cell[    3549] = 32'h0;  // 32'hcb0f1323;
    ram_cell[    3550] = 32'h0;  // 32'ha9838a12;
    ram_cell[    3551] = 32'h0;  // 32'hc3cdc6a5;
    ram_cell[    3552] = 32'h0;  // 32'h4ed5faf8;
    ram_cell[    3553] = 32'h0;  // 32'h2ffe48ea;
    ram_cell[    3554] = 32'h0;  // 32'h97c0015e;
    ram_cell[    3555] = 32'h0;  // 32'hc3af6722;
    ram_cell[    3556] = 32'h0;  // 32'hdddd4c50;
    ram_cell[    3557] = 32'h0;  // 32'h99d75286;
    ram_cell[    3558] = 32'h0;  // 32'hd7d5c211;
    ram_cell[    3559] = 32'h0;  // 32'h313c115f;
    ram_cell[    3560] = 32'h0;  // 32'he7d23463;
    ram_cell[    3561] = 32'h0;  // 32'h3cfce8cc;
    ram_cell[    3562] = 32'h0;  // 32'h292c6962;
    ram_cell[    3563] = 32'h0;  // 32'h41793288;
    ram_cell[    3564] = 32'h0;  // 32'hf2d2a50c;
    ram_cell[    3565] = 32'h0;  // 32'hc31af257;
    ram_cell[    3566] = 32'h0;  // 32'h882ca5e0;
    ram_cell[    3567] = 32'h0;  // 32'h6ab88de4;
    ram_cell[    3568] = 32'h0;  // 32'hc35c2b7f;
    ram_cell[    3569] = 32'h0;  // 32'hf79fae8b;
    ram_cell[    3570] = 32'h0;  // 32'h4330c6fe;
    ram_cell[    3571] = 32'h0;  // 32'h4c45f9f0;
    ram_cell[    3572] = 32'h0;  // 32'h3445172f;
    ram_cell[    3573] = 32'h0;  // 32'h91433504;
    ram_cell[    3574] = 32'h0;  // 32'ha36e3fb1;
    ram_cell[    3575] = 32'h0;  // 32'h32b7a89a;
    ram_cell[    3576] = 32'h0;  // 32'hc0f5bed3;
    ram_cell[    3577] = 32'h0;  // 32'h98f7f6db;
    ram_cell[    3578] = 32'h0;  // 32'ha567dd26;
    ram_cell[    3579] = 32'h0;  // 32'h6cc06e04;
    ram_cell[    3580] = 32'h0;  // 32'h3982da57;
    ram_cell[    3581] = 32'h0;  // 32'h6ec226f9;
    ram_cell[    3582] = 32'h0;  // 32'h2c739f0c;
    ram_cell[    3583] = 32'h0;  // 32'hec70a16b;
    ram_cell[    3584] = 32'h0;  // 32'ha156f4f0;
    ram_cell[    3585] = 32'h0;  // 32'hc11b5e1d;
    ram_cell[    3586] = 32'h0;  // 32'h9771425b;
    ram_cell[    3587] = 32'h0;  // 32'hd498f281;
    ram_cell[    3588] = 32'h0;  // 32'h13565e47;
    ram_cell[    3589] = 32'h0;  // 32'h985c9a31;
    ram_cell[    3590] = 32'h0;  // 32'h7e66071e;
    ram_cell[    3591] = 32'h0;  // 32'haaaf6167;
    ram_cell[    3592] = 32'h0;  // 32'hca3cc37f;
    ram_cell[    3593] = 32'h0;  // 32'h65c03ba8;
    ram_cell[    3594] = 32'h0;  // 32'h6b789a5d;
    ram_cell[    3595] = 32'h0;  // 32'hf88cb161;
    ram_cell[    3596] = 32'h0;  // 32'h182fafa9;
    ram_cell[    3597] = 32'h0;  // 32'h6f90cd2a;
    ram_cell[    3598] = 32'h0;  // 32'h34db2d44;
    ram_cell[    3599] = 32'h0;  // 32'habe3304a;
    ram_cell[    3600] = 32'h0;  // 32'h94dcbe17;
    ram_cell[    3601] = 32'h0;  // 32'h59e7c26b;
    ram_cell[    3602] = 32'h0;  // 32'h042453ad;
    ram_cell[    3603] = 32'h0;  // 32'h308b33cd;
    ram_cell[    3604] = 32'h0;  // 32'h909f2256;
    ram_cell[    3605] = 32'h0;  // 32'hcacab528;
    ram_cell[    3606] = 32'h0;  // 32'h5b6df67f;
    ram_cell[    3607] = 32'h0;  // 32'hf3694da1;
    ram_cell[    3608] = 32'h0;  // 32'h597c3521;
    ram_cell[    3609] = 32'h0;  // 32'h3c27f428;
    ram_cell[    3610] = 32'h0;  // 32'hdca7ef76;
    ram_cell[    3611] = 32'h0;  // 32'he67713ce;
    ram_cell[    3612] = 32'h0;  // 32'h106eccb6;
    ram_cell[    3613] = 32'h0;  // 32'h4be7dd5c;
    ram_cell[    3614] = 32'h0;  // 32'h2ca1bca9;
    ram_cell[    3615] = 32'h0;  // 32'ha7b2e39e;
    ram_cell[    3616] = 32'h0;  // 32'ha0532102;
    ram_cell[    3617] = 32'h0;  // 32'h1b7d3a4e;
    ram_cell[    3618] = 32'h0;  // 32'h5b0feaa8;
    ram_cell[    3619] = 32'h0;  // 32'hf32e5212;
    ram_cell[    3620] = 32'h0;  // 32'hb5cdeda5;
    ram_cell[    3621] = 32'h0;  // 32'hac91d163;
    ram_cell[    3622] = 32'h0;  // 32'hf0cb2009;
    ram_cell[    3623] = 32'h0;  // 32'h9202a9de;
    ram_cell[    3624] = 32'h0;  // 32'hd551e709;
    ram_cell[    3625] = 32'h0;  // 32'hf65185b0;
    ram_cell[    3626] = 32'h0;  // 32'h3cc81edb;
    ram_cell[    3627] = 32'h0;  // 32'h7dbfb8e2;
    ram_cell[    3628] = 32'h0;  // 32'h50d0160b;
    ram_cell[    3629] = 32'h0;  // 32'ha9897a31;
    ram_cell[    3630] = 32'h0;  // 32'h092c36e2;
    ram_cell[    3631] = 32'h0;  // 32'h3e60953e;
    ram_cell[    3632] = 32'h0;  // 32'hfef1a3a2;
    ram_cell[    3633] = 32'h0;  // 32'hda08be75;
    ram_cell[    3634] = 32'h0;  // 32'hfc45c45e;
    ram_cell[    3635] = 32'h0;  // 32'hff3b079c;
    ram_cell[    3636] = 32'h0;  // 32'h9bd941f4;
    ram_cell[    3637] = 32'h0;  // 32'hbed6ab83;
    ram_cell[    3638] = 32'h0;  // 32'h311bb451;
    ram_cell[    3639] = 32'h0;  // 32'h4d4d3ebd;
    ram_cell[    3640] = 32'h0;  // 32'h3b694a57;
    ram_cell[    3641] = 32'h0;  // 32'ha66ae74c;
    ram_cell[    3642] = 32'h0;  // 32'hcfca6334;
    ram_cell[    3643] = 32'h0;  // 32'h82239163;
    ram_cell[    3644] = 32'h0;  // 32'hc0fb77fe;
    ram_cell[    3645] = 32'h0;  // 32'h430783b4;
    ram_cell[    3646] = 32'h0;  // 32'h01aeb1cc;
    ram_cell[    3647] = 32'h0;  // 32'h262c70b2;
    ram_cell[    3648] = 32'h0;  // 32'hd14afc36;
    ram_cell[    3649] = 32'h0;  // 32'hf360ba79;
    ram_cell[    3650] = 32'h0;  // 32'h6647e50a;
    ram_cell[    3651] = 32'h0;  // 32'hfc639249;
    ram_cell[    3652] = 32'h0;  // 32'h091939f3;
    ram_cell[    3653] = 32'h0;  // 32'h36813445;
    ram_cell[    3654] = 32'h0;  // 32'he80fae33;
    ram_cell[    3655] = 32'h0;  // 32'h8c99312d;
    ram_cell[    3656] = 32'h0;  // 32'hda99f700;
    ram_cell[    3657] = 32'h0;  // 32'hd5ebea1e;
    ram_cell[    3658] = 32'h0;  // 32'hf86a45a3;
    ram_cell[    3659] = 32'h0;  // 32'hcf59ff25;
    ram_cell[    3660] = 32'h0;  // 32'h7b3a24f8;
    ram_cell[    3661] = 32'h0;  // 32'hc78af73e;
    ram_cell[    3662] = 32'h0;  // 32'he51f4965;
    ram_cell[    3663] = 32'h0;  // 32'h83e7aebb;
    ram_cell[    3664] = 32'h0;  // 32'h42ae5078;
    ram_cell[    3665] = 32'h0;  // 32'hac951840;
    ram_cell[    3666] = 32'h0;  // 32'ha61ff55c;
    ram_cell[    3667] = 32'h0;  // 32'h6379bbdc;
    ram_cell[    3668] = 32'h0;  // 32'h648eebd4;
    ram_cell[    3669] = 32'h0;  // 32'h3c55e531;
    ram_cell[    3670] = 32'h0;  // 32'h85f6e314;
    ram_cell[    3671] = 32'h0;  // 32'h48c843ee;
    ram_cell[    3672] = 32'h0;  // 32'h553ca3ce;
    ram_cell[    3673] = 32'h0;  // 32'hed902627;
    ram_cell[    3674] = 32'h0;  // 32'h41f78f92;
    ram_cell[    3675] = 32'h0;  // 32'h22f4523e;
    ram_cell[    3676] = 32'h0;  // 32'h49f78694;
    ram_cell[    3677] = 32'h0;  // 32'h9d791fcb;
    ram_cell[    3678] = 32'h0;  // 32'h38c6ce47;
    ram_cell[    3679] = 32'h0;  // 32'h60802ed3;
    ram_cell[    3680] = 32'h0;  // 32'ha6520920;
    ram_cell[    3681] = 32'h0;  // 32'he6c441ca;
    ram_cell[    3682] = 32'h0;  // 32'h3382faa3;
    ram_cell[    3683] = 32'h0;  // 32'had102098;
    ram_cell[    3684] = 32'h0;  // 32'h96bed9e2;
    ram_cell[    3685] = 32'h0;  // 32'hf2d66e20;
    ram_cell[    3686] = 32'h0;  // 32'h312559a4;
    ram_cell[    3687] = 32'h0;  // 32'h8d52a2d3;
    ram_cell[    3688] = 32'h0;  // 32'h835c832b;
    ram_cell[    3689] = 32'h0;  // 32'h5d559e09;
    ram_cell[    3690] = 32'h0;  // 32'h194dfcfe;
    ram_cell[    3691] = 32'h0;  // 32'ha7d22622;
    ram_cell[    3692] = 32'h0;  // 32'h49bf3803;
    ram_cell[    3693] = 32'h0;  // 32'h0544b067;
    ram_cell[    3694] = 32'h0;  // 32'h1645882b;
    ram_cell[    3695] = 32'h0;  // 32'h33526452;
    ram_cell[    3696] = 32'h0;  // 32'h9404f0da;
    ram_cell[    3697] = 32'h0;  // 32'hdeea43f2;
    ram_cell[    3698] = 32'h0;  // 32'h9d49c081;
    ram_cell[    3699] = 32'h0;  // 32'h4567cda5;
    ram_cell[    3700] = 32'h0;  // 32'h3309d3aa;
    ram_cell[    3701] = 32'h0;  // 32'hec59a967;
    ram_cell[    3702] = 32'h0;  // 32'hf7094fa4;
    ram_cell[    3703] = 32'h0;  // 32'h96a99708;
    ram_cell[    3704] = 32'h0;  // 32'ha4a00c7e;
    ram_cell[    3705] = 32'h0;  // 32'h8a35e770;
    ram_cell[    3706] = 32'h0;  // 32'h174e1e6a;
    ram_cell[    3707] = 32'h0;  // 32'h8063cf39;
    ram_cell[    3708] = 32'h0;  // 32'h2ac638b7;
    ram_cell[    3709] = 32'h0;  // 32'hf967877b;
    ram_cell[    3710] = 32'h0;  // 32'hdf088565;
    ram_cell[    3711] = 32'h0;  // 32'ha73eeb11;
    ram_cell[    3712] = 32'h0;  // 32'h71278c2b;
    ram_cell[    3713] = 32'h0;  // 32'h289d2c8d;
    ram_cell[    3714] = 32'h0;  // 32'h73800e6f;
    ram_cell[    3715] = 32'h0;  // 32'h0c880f02;
    ram_cell[    3716] = 32'h0;  // 32'ha686f849;
    ram_cell[    3717] = 32'h0;  // 32'h6fa82db8;
    ram_cell[    3718] = 32'h0;  // 32'h31df0e49;
    ram_cell[    3719] = 32'h0;  // 32'hc83b0fd1;
    ram_cell[    3720] = 32'h0;  // 32'h5d440817;
    ram_cell[    3721] = 32'h0;  // 32'h904787c3;
    ram_cell[    3722] = 32'h0;  // 32'h44f283f3;
    ram_cell[    3723] = 32'h0;  // 32'hd80adf90;
    ram_cell[    3724] = 32'h0;  // 32'h3bb79310;
    ram_cell[    3725] = 32'h0;  // 32'h75d03d57;
    ram_cell[    3726] = 32'h0;  // 32'hf1ac5afa;
    ram_cell[    3727] = 32'h0;  // 32'h123404ba;
    ram_cell[    3728] = 32'h0;  // 32'h6553a048;
    ram_cell[    3729] = 32'h0;  // 32'h46831f15;
    ram_cell[    3730] = 32'h0;  // 32'h70468480;
    ram_cell[    3731] = 32'h0;  // 32'hac39a609;
    ram_cell[    3732] = 32'h0;  // 32'h713b0994;
    ram_cell[    3733] = 32'h0;  // 32'ha15a1ce4;
    ram_cell[    3734] = 32'h0;  // 32'hff2ea10c;
    ram_cell[    3735] = 32'h0;  // 32'h0f40e86f;
    ram_cell[    3736] = 32'h0;  // 32'h9b8e611a;
    ram_cell[    3737] = 32'h0;  // 32'hed46aec2;
    ram_cell[    3738] = 32'h0;  // 32'h96d3deb9;
    ram_cell[    3739] = 32'h0;  // 32'h1da08dd8;
    ram_cell[    3740] = 32'h0;  // 32'hd40ef57d;
    ram_cell[    3741] = 32'h0;  // 32'h9c98bc0d;
    ram_cell[    3742] = 32'h0;  // 32'h64c1d604;
    ram_cell[    3743] = 32'h0;  // 32'h706e8ee1;
    ram_cell[    3744] = 32'h0;  // 32'h799c1d8c;
    ram_cell[    3745] = 32'h0;  // 32'h5a9fe9ef;
    ram_cell[    3746] = 32'h0;  // 32'h6ec5198c;
    ram_cell[    3747] = 32'h0;  // 32'hebceaa9d;
    ram_cell[    3748] = 32'h0;  // 32'ha8eabd50;
    ram_cell[    3749] = 32'h0;  // 32'h8e9f9904;
    ram_cell[    3750] = 32'h0;  // 32'h01917d38;
    ram_cell[    3751] = 32'h0;  // 32'h6e32fec9;
    ram_cell[    3752] = 32'h0;  // 32'h137a0c92;
    ram_cell[    3753] = 32'h0;  // 32'hff311c98;
    ram_cell[    3754] = 32'h0;  // 32'h5dbe9de1;
    ram_cell[    3755] = 32'h0;  // 32'he26b4068;
    ram_cell[    3756] = 32'h0;  // 32'hcd670a02;
    ram_cell[    3757] = 32'h0;  // 32'h018d6ed8;
    ram_cell[    3758] = 32'h0;  // 32'h25f0b46a;
    ram_cell[    3759] = 32'h0;  // 32'h2f1d839f;
    ram_cell[    3760] = 32'h0;  // 32'h293a356a;
    ram_cell[    3761] = 32'h0;  // 32'hd6825714;
    ram_cell[    3762] = 32'h0;  // 32'h179736c1;
    ram_cell[    3763] = 32'h0;  // 32'h96e03358;
    ram_cell[    3764] = 32'h0;  // 32'h2bf1d5d0;
    ram_cell[    3765] = 32'h0;  // 32'h373dc717;
    ram_cell[    3766] = 32'h0;  // 32'hd5721f29;
    ram_cell[    3767] = 32'h0;  // 32'h9ce0eb19;
    ram_cell[    3768] = 32'h0;  // 32'h84be51d7;
    ram_cell[    3769] = 32'h0;  // 32'h69d37a4f;
    ram_cell[    3770] = 32'h0;  // 32'h027f40d3;
    ram_cell[    3771] = 32'h0;  // 32'ha80324b1;
    ram_cell[    3772] = 32'h0;  // 32'he34eb0cf;
    ram_cell[    3773] = 32'h0;  // 32'h55004623;
    ram_cell[    3774] = 32'h0;  // 32'he0824ee2;
    ram_cell[    3775] = 32'h0;  // 32'h7ea02c16;
    ram_cell[    3776] = 32'h0;  // 32'hbe1d85d5;
    ram_cell[    3777] = 32'h0;  // 32'h09ffbe51;
    ram_cell[    3778] = 32'h0;  // 32'h4323a458;
    ram_cell[    3779] = 32'h0;  // 32'h80c68b70;
    ram_cell[    3780] = 32'h0;  // 32'hbcf8163a;
    ram_cell[    3781] = 32'h0;  // 32'h35bb62c5;
    ram_cell[    3782] = 32'h0;  // 32'h84604430;
    ram_cell[    3783] = 32'h0;  // 32'he36be259;
    ram_cell[    3784] = 32'h0;  // 32'hd5fbdb18;
    ram_cell[    3785] = 32'h0;  // 32'hfcdcc1de;
    ram_cell[    3786] = 32'h0;  // 32'hb0b99793;
    ram_cell[    3787] = 32'h0;  // 32'h4226ee57;
    ram_cell[    3788] = 32'h0;  // 32'h01c44bb4;
    ram_cell[    3789] = 32'h0;  // 32'h04054987;
    ram_cell[    3790] = 32'h0;  // 32'h9063a725;
    ram_cell[    3791] = 32'h0;  // 32'h4efa383e;
    ram_cell[    3792] = 32'h0;  // 32'ha667f1ad;
    ram_cell[    3793] = 32'h0;  // 32'h38577866;
    ram_cell[    3794] = 32'h0;  // 32'he0c77194;
    ram_cell[    3795] = 32'h0;  // 32'h6eb52760;
    ram_cell[    3796] = 32'h0;  // 32'haa0e3206;
    ram_cell[    3797] = 32'h0;  // 32'hcb641ff5;
    ram_cell[    3798] = 32'h0;  // 32'h16793c12;
    ram_cell[    3799] = 32'h0;  // 32'hb187dd32;
    ram_cell[    3800] = 32'h0;  // 32'h4ebaf544;
    ram_cell[    3801] = 32'h0;  // 32'h724b3274;
    ram_cell[    3802] = 32'h0;  // 32'he4f0a2d3;
    ram_cell[    3803] = 32'h0;  // 32'h776c0487;
    ram_cell[    3804] = 32'h0;  // 32'h80779127;
    ram_cell[    3805] = 32'h0;  // 32'ha0c6d9ad;
    ram_cell[    3806] = 32'h0;  // 32'h48aef833;
    ram_cell[    3807] = 32'h0;  // 32'hf59fdb83;
    ram_cell[    3808] = 32'h0;  // 32'h72b56eac;
    ram_cell[    3809] = 32'h0;  // 32'h48f47b98;
    ram_cell[    3810] = 32'h0;  // 32'hc00f5b87;
    ram_cell[    3811] = 32'h0;  // 32'h6ef59600;
    ram_cell[    3812] = 32'h0;  // 32'h9ad2c608;
    ram_cell[    3813] = 32'h0;  // 32'h7929e9e6;
    ram_cell[    3814] = 32'h0;  // 32'h35b297a6;
    ram_cell[    3815] = 32'h0;  // 32'h6e489ad0;
    ram_cell[    3816] = 32'h0;  // 32'hf8b2fba1;
    ram_cell[    3817] = 32'h0;  // 32'hbea37976;
    ram_cell[    3818] = 32'h0;  // 32'h4fa55da9;
    ram_cell[    3819] = 32'h0;  // 32'ha38fa5fc;
    ram_cell[    3820] = 32'h0;  // 32'hbe49ebe7;
    ram_cell[    3821] = 32'h0;  // 32'h2dbdebc0;
    ram_cell[    3822] = 32'h0;  // 32'h093e75d3;
    ram_cell[    3823] = 32'h0;  // 32'h90248f95;
    ram_cell[    3824] = 32'h0;  // 32'hf576e11b;
    ram_cell[    3825] = 32'h0;  // 32'he1687d95;
    ram_cell[    3826] = 32'h0;  // 32'hf9e3a457;
    ram_cell[    3827] = 32'h0;  // 32'h1042daf3;
    ram_cell[    3828] = 32'h0;  // 32'hbb00c88e;
    ram_cell[    3829] = 32'h0;  // 32'h6c50eeee;
    ram_cell[    3830] = 32'h0;  // 32'h8152ec7a;
    ram_cell[    3831] = 32'h0;  // 32'h7419a313;
    ram_cell[    3832] = 32'h0;  // 32'hb93f6db2;
    ram_cell[    3833] = 32'h0;  // 32'h08cb7534;
    ram_cell[    3834] = 32'h0;  // 32'h1134930e;
    ram_cell[    3835] = 32'h0;  // 32'h1057f64f;
    ram_cell[    3836] = 32'h0;  // 32'hf9607025;
    ram_cell[    3837] = 32'h0;  // 32'h393ade55;
    ram_cell[    3838] = 32'h0;  // 32'h31c2a6de;
    ram_cell[    3839] = 32'h0;  // 32'h9237f7d4;
    ram_cell[    3840] = 32'h0;  // 32'heee67f17;
    ram_cell[    3841] = 32'h0;  // 32'h105bc882;
    ram_cell[    3842] = 32'h0;  // 32'hcf18cac1;
    ram_cell[    3843] = 32'h0;  // 32'he592c788;
    ram_cell[    3844] = 32'h0;  // 32'h31989a7c;
    ram_cell[    3845] = 32'h0;  // 32'h6b229bee;
    ram_cell[    3846] = 32'h0;  // 32'h6df036ab;
    ram_cell[    3847] = 32'h0;  // 32'h1603d721;
    ram_cell[    3848] = 32'h0;  // 32'heead1137;
    ram_cell[    3849] = 32'h0;  // 32'he4021a39;
    ram_cell[    3850] = 32'h0;  // 32'hfaed5ef4;
    ram_cell[    3851] = 32'h0;  // 32'h794aaa5e;
    ram_cell[    3852] = 32'h0;  // 32'h05c20601;
    ram_cell[    3853] = 32'h0;  // 32'hde2c8cb6;
    ram_cell[    3854] = 32'h0;  // 32'h5deb6bd7;
    ram_cell[    3855] = 32'h0;  // 32'haad5fee8;
    ram_cell[    3856] = 32'h0;  // 32'h7a02d622;
    ram_cell[    3857] = 32'h0;  // 32'hda8c684b;
    ram_cell[    3858] = 32'h0;  // 32'h4f2fd8db;
    ram_cell[    3859] = 32'h0;  // 32'hf484fc68;
    ram_cell[    3860] = 32'h0;  // 32'h9e7d83d4;
    ram_cell[    3861] = 32'h0;  // 32'hbe774e7a;
    ram_cell[    3862] = 32'h0;  // 32'hac5667ab;
    ram_cell[    3863] = 32'h0;  // 32'h2386d957;
    ram_cell[    3864] = 32'h0;  // 32'hd516fea5;
    ram_cell[    3865] = 32'h0;  // 32'h77a557c4;
    ram_cell[    3866] = 32'h0;  // 32'h3bf069ff;
    ram_cell[    3867] = 32'h0;  // 32'hf17f6f15;
    ram_cell[    3868] = 32'h0;  // 32'ha4b9380c;
    ram_cell[    3869] = 32'h0;  // 32'h89c0add4;
    ram_cell[    3870] = 32'h0;  // 32'h97b40365;
    ram_cell[    3871] = 32'h0;  // 32'h0a8ec99c;
    ram_cell[    3872] = 32'h0;  // 32'hf799031e;
    ram_cell[    3873] = 32'h0;  // 32'he399e92a;
    ram_cell[    3874] = 32'h0;  // 32'h5fb00811;
    ram_cell[    3875] = 32'h0;  // 32'h6363dcf2;
    ram_cell[    3876] = 32'h0;  // 32'h852c2e74;
    ram_cell[    3877] = 32'h0;  // 32'h7f376690;
    ram_cell[    3878] = 32'h0;  // 32'hc1b38b34;
    ram_cell[    3879] = 32'h0;  // 32'h661cbdad;
    ram_cell[    3880] = 32'h0;  // 32'h30a7dd7f;
    ram_cell[    3881] = 32'h0;  // 32'h421bd4c6;
    ram_cell[    3882] = 32'h0;  // 32'hd7655a3e;
    ram_cell[    3883] = 32'h0;  // 32'had9c99d1;
    ram_cell[    3884] = 32'h0;  // 32'h13502d32;
    ram_cell[    3885] = 32'h0;  // 32'h20910853;
    ram_cell[    3886] = 32'h0;  // 32'h64e4eb3d;
    ram_cell[    3887] = 32'h0;  // 32'he1d0ca6e;
    ram_cell[    3888] = 32'h0;  // 32'h0652fb0c;
    ram_cell[    3889] = 32'h0;  // 32'h600b96d6;
    ram_cell[    3890] = 32'h0;  // 32'h6a6bc91d;
    ram_cell[    3891] = 32'h0;  // 32'hfeaf0a41;
    ram_cell[    3892] = 32'h0;  // 32'h58160714;
    ram_cell[    3893] = 32'h0;  // 32'h5bf6c5aa;
    ram_cell[    3894] = 32'h0;  // 32'heccd9899;
    ram_cell[    3895] = 32'h0;  // 32'h4447dd23;
    ram_cell[    3896] = 32'h0;  // 32'h5c3e1354;
    ram_cell[    3897] = 32'h0;  // 32'h13983e91;
    ram_cell[    3898] = 32'h0;  // 32'h29e7b561;
    ram_cell[    3899] = 32'h0;  // 32'h143de51a;
    ram_cell[    3900] = 32'h0;  // 32'hd2ddb729;
    ram_cell[    3901] = 32'h0;  // 32'h6cbf64cf;
    ram_cell[    3902] = 32'h0;  // 32'h3b461625;
    ram_cell[    3903] = 32'h0;  // 32'hc225d7f3;
    ram_cell[    3904] = 32'h0;  // 32'h0c60c682;
    ram_cell[    3905] = 32'h0;  // 32'h6d560e4b;
    ram_cell[    3906] = 32'h0;  // 32'h5b17e7ae;
    ram_cell[    3907] = 32'h0;  // 32'h533b6778;
    ram_cell[    3908] = 32'h0;  // 32'hd804ae46;
    ram_cell[    3909] = 32'h0;  // 32'hdf59edfb;
    ram_cell[    3910] = 32'h0;  // 32'h072820f1;
    ram_cell[    3911] = 32'h0;  // 32'h8e21f5c0;
    ram_cell[    3912] = 32'h0;  // 32'hfea7ab42;
    ram_cell[    3913] = 32'h0;  // 32'h4be47732;
    ram_cell[    3914] = 32'h0;  // 32'h7aa8bc3c;
    ram_cell[    3915] = 32'h0;  // 32'h746e971c;
    ram_cell[    3916] = 32'h0;  // 32'h4d88c2c0;
    ram_cell[    3917] = 32'h0;  // 32'h75216c92;
    ram_cell[    3918] = 32'h0;  // 32'h9ba523d4;
    ram_cell[    3919] = 32'h0;  // 32'h5ed5365b;
    ram_cell[    3920] = 32'h0;  // 32'hf36a7bc6;
    ram_cell[    3921] = 32'h0;  // 32'h87dc4fcf;
    ram_cell[    3922] = 32'h0;  // 32'h3c18b3a2;
    ram_cell[    3923] = 32'h0;  // 32'h5aa567bc;
    ram_cell[    3924] = 32'h0;  // 32'h9faa77c8;
    ram_cell[    3925] = 32'h0;  // 32'hb0e4917c;
    ram_cell[    3926] = 32'h0;  // 32'h6984cceb;
    ram_cell[    3927] = 32'h0;  // 32'h4eece4de;
    ram_cell[    3928] = 32'h0;  // 32'hde8bac2c;
    ram_cell[    3929] = 32'h0;  // 32'hb9aa7ab5;
    ram_cell[    3930] = 32'h0;  // 32'h2feef30c;
    ram_cell[    3931] = 32'h0;  // 32'hd29b5775;
    ram_cell[    3932] = 32'h0;  // 32'he17f85b2;
    ram_cell[    3933] = 32'h0;  // 32'he90d61c2;
    ram_cell[    3934] = 32'h0;  // 32'h3566b3ca;
    ram_cell[    3935] = 32'h0;  // 32'h5ef6e0c7;
    ram_cell[    3936] = 32'h0;  // 32'he4bf5f7d;
    ram_cell[    3937] = 32'h0;  // 32'hf0c39fd0;
    ram_cell[    3938] = 32'h0;  // 32'h40848ccb;
    ram_cell[    3939] = 32'h0;  // 32'h48910679;
    ram_cell[    3940] = 32'h0;  // 32'h74d6682d;
    ram_cell[    3941] = 32'h0;  // 32'h3af0ce7f;
    ram_cell[    3942] = 32'h0;  // 32'hcb171c90;
    ram_cell[    3943] = 32'h0;  // 32'h012b079a;
    ram_cell[    3944] = 32'h0;  // 32'h1cd3bcdc;
    ram_cell[    3945] = 32'h0;  // 32'h3a036645;
    ram_cell[    3946] = 32'h0;  // 32'h8b560234;
    ram_cell[    3947] = 32'h0;  // 32'hd9c9c497;
    ram_cell[    3948] = 32'h0;  // 32'h193f0334;
    ram_cell[    3949] = 32'h0;  // 32'h3d98cc31;
    ram_cell[    3950] = 32'h0;  // 32'hddc9e2ae;
    ram_cell[    3951] = 32'h0;  // 32'hb3fe8091;
    ram_cell[    3952] = 32'h0;  // 32'had0565f5;
    ram_cell[    3953] = 32'h0;  // 32'hfca82d56;
    ram_cell[    3954] = 32'h0;  // 32'hc0c674fb;
    ram_cell[    3955] = 32'h0;  // 32'h5a39d131;
    ram_cell[    3956] = 32'h0;  // 32'h4fd096e3;
    ram_cell[    3957] = 32'h0;  // 32'h0bc016df;
    ram_cell[    3958] = 32'h0;  // 32'h75b3f118;
    ram_cell[    3959] = 32'h0;  // 32'h26498b66;
    ram_cell[    3960] = 32'h0;  // 32'hf2813114;
    ram_cell[    3961] = 32'h0;  // 32'h57c6682a;
    ram_cell[    3962] = 32'h0;  // 32'h1fb2d202;
    ram_cell[    3963] = 32'h0;  // 32'h8385190c;
    ram_cell[    3964] = 32'h0;  // 32'h18a6bc01;
    ram_cell[    3965] = 32'h0;  // 32'h8dbc1d92;
    ram_cell[    3966] = 32'h0;  // 32'he34dab29;
    ram_cell[    3967] = 32'h0;  // 32'hab675476;
    ram_cell[    3968] = 32'h0;  // 32'hb55bb94f;
    ram_cell[    3969] = 32'h0;  // 32'hfee8544b;
    ram_cell[    3970] = 32'h0;  // 32'h54cae477;
    ram_cell[    3971] = 32'h0;  // 32'hf1b76aad;
    ram_cell[    3972] = 32'h0;  // 32'hf63a33bf;
    ram_cell[    3973] = 32'h0;  // 32'h155e9939;
    ram_cell[    3974] = 32'h0;  // 32'hea07ad0e;
    ram_cell[    3975] = 32'h0;  // 32'h7407d519;
    ram_cell[    3976] = 32'h0;  // 32'h17c44927;
    ram_cell[    3977] = 32'h0;  // 32'h6f237069;
    ram_cell[    3978] = 32'h0;  // 32'h4a6218ea;
    ram_cell[    3979] = 32'h0;  // 32'h39b95218;
    ram_cell[    3980] = 32'h0;  // 32'h6e392b59;
    ram_cell[    3981] = 32'h0;  // 32'ha3fb1f6f;
    ram_cell[    3982] = 32'h0;  // 32'h54973a86;
    ram_cell[    3983] = 32'h0;  // 32'h83b61082;
    ram_cell[    3984] = 32'h0;  // 32'h64a7247f;
    ram_cell[    3985] = 32'h0;  // 32'h0f3d5968;
    ram_cell[    3986] = 32'h0;  // 32'hea2081e4;
    ram_cell[    3987] = 32'h0;  // 32'h054e01a1;
    ram_cell[    3988] = 32'h0;  // 32'haa3e0fe0;
    ram_cell[    3989] = 32'h0;  // 32'h8e3b660e;
    ram_cell[    3990] = 32'h0;  // 32'hea5405a3;
    ram_cell[    3991] = 32'h0;  // 32'hf2ec639d;
    ram_cell[    3992] = 32'h0;  // 32'h3c76d1ea;
    ram_cell[    3993] = 32'h0;  // 32'hdfeaa567;
    ram_cell[    3994] = 32'h0;  // 32'ha2c4ac63;
    ram_cell[    3995] = 32'h0;  // 32'h84b54790;
    ram_cell[    3996] = 32'h0;  // 32'h82f93a48;
    ram_cell[    3997] = 32'h0;  // 32'hb1593802;
    ram_cell[    3998] = 32'h0;  // 32'hb4d0cf05;
    ram_cell[    3999] = 32'h0;  // 32'h7c13984e;
    ram_cell[    4000] = 32'h0;  // 32'h38efa3a7;
    ram_cell[    4001] = 32'h0;  // 32'h162dba8f;
    ram_cell[    4002] = 32'h0;  // 32'h835b4c02;
    ram_cell[    4003] = 32'h0;  // 32'h3eecb80f;
    ram_cell[    4004] = 32'h0;  // 32'hbd2e1727;
    ram_cell[    4005] = 32'h0;  // 32'h9986b1d5;
    ram_cell[    4006] = 32'h0;  // 32'h01c39cef;
    ram_cell[    4007] = 32'h0;  // 32'hc671d2ce;
    ram_cell[    4008] = 32'h0;  // 32'h0b9737d2;
    ram_cell[    4009] = 32'h0;  // 32'hca00f8a2;
    ram_cell[    4010] = 32'h0;  // 32'hc1775347;
    ram_cell[    4011] = 32'h0;  // 32'hd2bd1892;
    ram_cell[    4012] = 32'h0;  // 32'hf67d7fdb;
    ram_cell[    4013] = 32'h0;  // 32'hc1c40b94;
    ram_cell[    4014] = 32'h0;  // 32'hea76e4a0;
    ram_cell[    4015] = 32'h0;  // 32'hdbf46b4e;
    ram_cell[    4016] = 32'h0;  // 32'h642e85fa;
    ram_cell[    4017] = 32'h0;  // 32'haebed146;
    ram_cell[    4018] = 32'h0;  // 32'hbb214ff1;
    ram_cell[    4019] = 32'h0;  // 32'hfcf00537;
    ram_cell[    4020] = 32'h0;  // 32'h870fa6a5;
    ram_cell[    4021] = 32'h0;  // 32'h0d44aa3d;
    ram_cell[    4022] = 32'h0;  // 32'hf4dab4a2;
    ram_cell[    4023] = 32'h0;  // 32'hb5eca3a1;
    ram_cell[    4024] = 32'h0;  // 32'h1a8ffa73;
    ram_cell[    4025] = 32'h0;  // 32'h1f30c0ae;
    ram_cell[    4026] = 32'h0;  // 32'hd4127c98;
    ram_cell[    4027] = 32'h0;  // 32'h1bb41fe5;
    ram_cell[    4028] = 32'h0;  // 32'hc88333bb;
    ram_cell[    4029] = 32'h0;  // 32'hc7683a87;
    ram_cell[    4030] = 32'h0;  // 32'h8c024c1f;
    ram_cell[    4031] = 32'h0;  // 32'h85b61e1d;
    ram_cell[    4032] = 32'h0;  // 32'h9aa6f31e;
    ram_cell[    4033] = 32'h0;  // 32'hc76d71b0;
    ram_cell[    4034] = 32'h0;  // 32'h2a5fb788;
    ram_cell[    4035] = 32'h0;  // 32'h4e079e57;
    ram_cell[    4036] = 32'h0;  // 32'hf0dec1fa;
    ram_cell[    4037] = 32'h0;  // 32'hbaf3f854;
    ram_cell[    4038] = 32'h0;  // 32'h3b8e6a98;
    ram_cell[    4039] = 32'h0;  // 32'hbf646dc6;
    ram_cell[    4040] = 32'h0;  // 32'hbc80f35b;
    ram_cell[    4041] = 32'h0;  // 32'h9e6bd3b5;
    ram_cell[    4042] = 32'h0;  // 32'hd6d4361f;
    ram_cell[    4043] = 32'h0;  // 32'ha013ccac;
    ram_cell[    4044] = 32'h0;  // 32'ha508ad81;
    ram_cell[    4045] = 32'h0;  // 32'h3554847d;
    ram_cell[    4046] = 32'h0;  // 32'h538a80ce;
    ram_cell[    4047] = 32'h0;  // 32'h91e9dbf4;
    ram_cell[    4048] = 32'h0;  // 32'hbf413d8d;
    ram_cell[    4049] = 32'h0;  // 32'he81bb27a;
    ram_cell[    4050] = 32'h0;  // 32'h3cf89c32;
    ram_cell[    4051] = 32'h0;  // 32'h83790016;
    ram_cell[    4052] = 32'h0;  // 32'h753a8ae4;
    ram_cell[    4053] = 32'h0;  // 32'h5dc899e0;
    ram_cell[    4054] = 32'h0;  // 32'hf9333ac9;
    ram_cell[    4055] = 32'h0;  // 32'hfb91e7ba;
    ram_cell[    4056] = 32'h0;  // 32'hdcf77d20;
    ram_cell[    4057] = 32'h0;  // 32'h3e918147;
    ram_cell[    4058] = 32'h0;  // 32'h10045865;
    ram_cell[    4059] = 32'h0;  // 32'h61f3c227;
    ram_cell[    4060] = 32'h0;  // 32'ha7f6b0e5;
    ram_cell[    4061] = 32'h0;  // 32'h1b301f61;
    ram_cell[    4062] = 32'h0;  // 32'hc0c9af74;
    ram_cell[    4063] = 32'h0;  // 32'h089c9c98;
    ram_cell[    4064] = 32'h0;  // 32'h8c30c573;
    ram_cell[    4065] = 32'h0;  // 32'h57c16878;
    ram_cell[    4066] = 32'h0;  // 32'h6aa8d494;
    ram_cell[    4067] = 32'h0;  // 32'h9e08ab6b;
    ram_cell[    4068] = 32'h0;  // 32'hea941907;
    ram_cell[    4069] = 32'h0;  // 32'h177ae740;
    ram_cell[    4070] = 32'h0;  // 32'hd03b144e;
    ram_cell[    4071] = 32'h0;  // 32'h1fb84c31;
    ram_cell[    4072] = 32'h0;  // 32'h4c74bcc3;
    ram_cell[    4073] = 32'h0;  // 32'h39a0e60a;
    ram_cell[    4074] = 32'h0;  // 32'hf423ca90;
    ram_cell[    4075] = 32'h0;  // 32'he0d9a5e2;
    ram_cell[    4076] = 32'h0;  // 32'h405b0a84;
    ram_cell[    4077] = 32'h0;  // 32'h767284ca;
    ram_cell[    4078] = 32'h0;  // 32'h0d96f271;
    ram_cell[    4079] = 32'h0;  // 32'h9e74983e;
    ram_cell[    4080] = 32'h0;  // 32'h9209e19a;
    ram_cell[    4081] = 32'h0;  // 32'h0ed4afa3;
    ram_cell[    4082] = 32'h0;  // 32'h4be227d0;
    ram_cell[    4083] = 32'h0;  // 32'h4040f658;
    ram_cell[    4084] = 32'h0;  // 32'h3a6269be;
    ram_cell[    4085] = 32'h0;  // 32'hf33804ab;
    ram_cell[    4086] = 32'h0;  // 32'hb94eee96;
    ram_cell[    4087] = 32'h0;  // 32'h90f98d0f;
    ram_cell[    4088] = 32'h0;  // 32'h7ede4eba;
    ram_cell[    4089] = 32'h0;  // 32'he51b0d9f;
    ram_cell[    4090] = 32'h0;  // 32'h51bc1e49;
    ram_cell[    4091] = 32'h0;  // 32'h145ccac5;
    ram_cell[    4092] = 32'h0;  // 32'h357e75a8;
    ram_cell[    4093] = 32'h0;  // 32'h5c5fb567;
    ram_cell[    4094] = 32'h0;  // 32'h18bc9d52;
    ram_cell[    4095] = 32'h0;  // 32'h8994b6db;
    // src matrix A
    ram_cell[    4096] = 32'ha932470e;
    ram_cell[    4097] = 32'h1989cff9;
    ram_cell[    4098] = 32'hf2e6f37f;
    ram_cell[    4099] = 32'h67d9f400;
    ram_cell[    4100] = 32'hb989c3d5;
    ram_cell[    4101] = 32'h2aea0015;
    ram_cell[    4102] = 32'h5faec516;
    ram_cell[    4103] = 32'h6c4a5e86;
    ram_cell[    4104] = 32'h7b4039ac;
    ram_cell[    4105] = 32'h23229782;
    ram_cell[    4106] = 32'hd882d71a;
    ram_cell[    4107] = 32'hdb3ff17d;
    ram_cell[    4108] = 32'ha1b12c5f;
    ram_cell[    4109] = 32'ha0dbdcea;
    ram_cell[    4110] = 32'h160725c5;
    ram_cell[    4111] = 32'hfdfec3ba;
    ram_cell[    4112] = 32'heac7045b;
    ram_cell[    4113] = 32'h38fb6dfc;
    ram_cell[    4114] = 32'haff29321;
    ram_cell[    4115] = 32'h4604b780;
    ram_cell[    4116] = 32'hd11b010b;
    ram_cell[    4117] = 32'h3f0c99b4;
    ram_cell[    4118] = 32'hbd32a926;
    ram_cell[    4119] = 32'h5ee3e375;
    ram_cell[    4120] = 32'h5afcd49c;
    ram_cell[    4121] = 32'hbb3e022a;
    ram_cell[    4122] = 32'h19de444f;
    ram_cell[    4123] = 32'h12512d26;
    ram_cell[    4124] = 32'h45ded948;
    ram_cell[    4125] = 32'h9f66071b;
    ram_cell[    4126] = 32'h119d104a;
    ram_cell[    4127] = 32'h1324a047;
    ram_cell[    4128] = 32'hc0d540f6;
    ram_cell[    4129] = 32'h9d4aa704;
    ram_cell[    4130] = 32'h1eb15df7;
    ram_cell[    4131] = 32'hd5cf5d99;
    ram_cell[    4132] = 32'h82de508d;
    ram_cell[    4133] = 32'h40b0f519;
    ram_cell[    4134] = 32'hbbb9120c;
    ram_cell[    4135] = 32'h6f42c9b2;
    ram_cell[    4136] = 32'h58d41c7e;
    ram_cell[    4137] = 32'hf05ee1da;
    ram_cell[    4138] = 32'h1dccbebc;
    ram_cell[    4139] = 32'hb7122261;
    ram_cell[    4140] = 32'h01c08c3d;
    ram_cell[    4141] = 32'h2340221e;
    ram_cell[    4142] = 32'h0e1673ce;
    ram_cell[    4143] = 32'h250886bd;
    ram_cell[    4144] = 32'hf8dacbc6;
    ram_cell[    4145] = 32'h128557d0;
    ram_cell[    4146] = 32'h76a02048;
    ram_cell[    4147] = 32'h30d54fae;
    ram_cell[    4148] = 32'hfa96a628;
    ram_cell[    4149] = 32'h210b9cc2;
    ram_cell[    4150] = 32'hf58635b0;
    ram_cell[    4151] = 32'hc1e6fcf2;
    ram_cell[    4152] = 32'hcadb7a67;
    ram_cell[    4153] = 32'h48ba1af4;
    ram_cell[    4154] = 32'h5caa95f2;
    ram_cell[    4155] = 32'habb292d8;
    ram_cell[    4156] = 32'h46ade337;
    ram_cell[    4157] = 32'h6dedf511;
    ram_cell[    4158] = 32'hcce22e0f;
    ram_cell[    4159] = 32'h5650f4c4;
    ram_cell[    4160] = 32'h7624cd95;
    ram_cell[    4161] = 32'h466407f1;
    ram_cell[    4162] = 32'h2e08e0d7;
    ram_cell[    4163] = 32'hd2a5b7dd;
    ram_cell[    4164] = 32'h333f899c;
    ram_cell[    4165] = 32'h9f4a3c6f;
    ram_cell[    4166] = 32'h886aac2a;
    ram_cell[    4167] = 32'hd7c0341d;
    ram_cell[    4168] = 32'h2b92edb7;
    ram_cell[    4169] = 32'hdcb8a34b;
    ram_cell[    4170] = 32'h3e184694;
    ram_cell[    4171] = 32'h78c3a098;
    ram_cell[    4172] = 32'hd8df35b6;
    ram_cell[    4173] = 32'h9d4b0aae;
    ram_cell[    4174] = 32'hb1271e87;
    ram_cell[    4175] = 32'h7d15c73a;
    ram_cell[    4176] = 32'h0fc6d7a5;
    ram_cell[    4177] = 32'hfa9c663c;
    ram_cell[    4178] = 32'hf3aa118c;
    ram_cell[    4179] = 32'hbbe76ca8;
    ram_cell[    4180] = 32'hbdace662;
    ram_cell[    4181] = 32'hbd30a026;
    ram_cell[    4182] = 32'h9b1a8969;
    ram_cell[    4183] = 32'h3a7d9bb4;
    ram_cell[    4184] = 32'hb0f90a5b;
    ram_cell[    4185] = 32'hb451208c;
    ram_cell[    4186] = 32'h735db2fa;
    ram_cell[    4187] = 32'hf1fbb749;
    ram_cell[    4188] = 32'hb219dc15;
    ram_cell[    4189] = 32'hafdf0c0e;
    ram_cell[    4190] = 32'h22b4df14;
    ram_cell[    4191] = 32'h5e829edb;
    ram_cell[    4192] = 32'h48657a6a;
    ram_cell[    4193] = 32'h9ca653f0;
    ram_cell[    4194] = 32'hdd638351;
    ram_cell[    4195] = 32'h711c814b;
    ram_cell[    4196] = 32'h797bb9b5;
    ram_cell[    4197] = 32'hcc251738;
    ram_cell[    4198] = 32'he44b4c2b;
    ram_cell[    4199] = 32'h4d953907;
    ram_cell[    4200] = 32'hf9d5b801;
    ram_cell[    4201] = 32'ha8e0dd1e;
    ram_cell[    4202] = 32'h1dc5e09e;
    ram_cell[    4203] = 32'h0323edcf;
    ram_cell[    4204] = 32'h2afde993;
    ram_cell[    4205] = 32'he19d07a2;
    ram_cell[    4206] = 32'hcd9e0d39;
    ram_cell[    4207] = 32'hba313d10;
    ram_cell[    4208] = 32'hd6318bcb;
    ram_cell[    4209] = 32'hc24beb00;
    ram_cell[    4210] = 32'hceb34235;
    ram_cell[    4211] = 32'ha09ec97a;
    ram_cell[    4212] = 32'hed6021b6;
    ram_cell[    4213] = 32'h16a51a81;
    ram_cell[    4214] = 32'hf55ea389;
    ram_cell[    4215] = 32'h85d49677;
    ram_cell[    4216] = 32'heafdb1e0;
    ram_cell[    4217] = 32'h5f6c4588;
    ram_cell[    4218] = 32'h5cb38bbc;
    ram_cell[    4219] = 32'h4fa90448;
    ram_cell[    4220] = 32'hc32257e5;
    ram_cell[    4221] = 32'h4e65d5e3;
    ram_cell[    4222] = 32'haa8a2509;
    ram_cell[    4223] = 32'h6b5a21d3;
    ram_cell[    4224] = 32'h89983ac0;
    ram_cell[    4225] = 32'h68f87512;
    ram_cell[    4226] = 32'h41949a08;
    ram_cell[    4227] = 32'hca51e405;
    ram_cell[    4228] = 32'h0dd488fc;
    ram_cell[    4229] = 32'he24c4ba0;
    ram_cell[    4230] = 32'hc1e13ef8;
    ram_cell[    4231] = 32'h39a4b62a;
    ram_cell[    4232] = 32'h65387ea9;
    ram_cell[    4233] = 32'h5e45aaa3;
    ram_cell[    4234] = 32'h124f8e81;
    ram_cell[    4235] = 32'h47242ee2;
    ram_cell[    4236] = 32'h2ed80ced;
    ram_cell[    4237] = 32'h19f4aa81;
    ram_cell[    4238] = 32'h96f48cf9;
    ram_cell[    4239] = 32'h1147dc71;
    ram_cell[    4240] = 32'hbbd4deda;
    ram_cell[    4241] = 32'hfa98ef3c;
    ram_cell[    4242] = 32'hdac6e924;
    ram_cell[    4243] = 32'hf9be2149;
    ram_cell[    4244] = 32'h6a442078;
    ram_cell[    4245] = 32'h2f5138b5;
    ram_cell[    4246] = 32'h926dd394;
    ram_cell[    4247] = 32'h6c1fa154;
    ram_cell[    4248] = 32'hd68fa95f;
    ram_cell[    4249] = 32'hd16b1954;
    ram_cell[    4250] = 32'h15e2a08f;
    ram_cell[    4251] = 32'h8d047cdc;
    ram_cell[    4252] = 32'h4bad57e7;
    ram_cell[    4253] = 32'h500493f6;
    ram_cell[    4254] = 32'h737f12e9;
    ram_cell[    4255] = 32'h2b6a7bae;
    ram_cell[    4256] = 32'h16b1d82e;
    ram_cell[    4257] = 32'h9e6371de;
    ram_cell[    4258] = 32'hcbe235a5;
    ram_cell[    4259] = 32'h859f19e6;
    ram_cell[    4260] = 32'hb5475238;
    ram_cell[    4261] = 32'hb707466e;
    ram_cell[    4262] = 32'h108168e3;
    ram_cell[    4263] = 32'hdd37fe90;
    ram_cell[    4264] = 32'h0eff798a;
    ram_cell[    4265] = 32'h19209342;
    ram_cell[    4266] = 32'h9d649747;
    ram_cell[    4267] = 32'h9a52d81f;
    ram_cell[    4268] = 32'h0a11a091;
    ram_cell[    4269] = 32'hccc4ab7b;
    ram_cell[    4270] = 32'h954794b0;
    ram_cell[    4271] = 32'hd6bf3e47;
    ram_cell[    4272] = 32'h29af0267;
    ram_cell[    4273] = 32'hf3943e18;
    ram_cell[    4274] = 32'h76ab6e36;
    ram_cell[    4275] = 32'h92f2522e;
    ram_cell[    4276] = 32'h3105aeea;
    ram_cell[    4277] = 32'hed536bae;
    ram_cell[    4278] = 32'h5874a5e6;
    ram_cell[    4279] = 32'h8387e983;
    ram_cell[    4280] = 32'h694d1990;
    ram_cell[    4281] = 32'hc60165ba;
    ram_cell[    4282] = 32'h1eb20253;
    ram_cell[    4283] = 32'h2b0382dd;
    ram_cell[    4284] = 32'hf92529b8;
    ram_cell[    4285] = 32'he0fea797;
    ram_cell[    4286] = 32'h4ee5baf9;
    ram_cell[    4287] = 32'ha525a7f3;
    ram_cell[    4288] = 32'h2b7aa3db;
    ram_cell[    4289] = 32'h769c36d0;
    ram_cell[    4290] = 32'h806a2458;
    ram_cell[    4291] = 32'h951a60ab;
    ram_cell[    4292] = 32'hc24a4bd8;
    ram_cell[    4293] = 32'ha2af7ea6;
    ram_cell[    4294] = 32'h9b9cf0fd;
    ram_cell[    4295] = 32'he01e5ee6;
    ram_cell[    4296] = 32'h04df8b2f;
    ram_cell[    4297] = 32'h14de8679;
    ram_cell[    4298] = 32'hf69a7cdd;
    ram_cell[    4299] = 32'h13cfeafe;
    ram_cell[    4300] = 32'h24e46faa;
    ram_cell[    4301] = 32'h24f2afb7;
    ram_cell[    4302] = 32'h7593b002;
    ram_cell[    4303] = 32'hc65602e4;
    ram_cell[    4304] = 32'h5ee71831;
    ram_cell[    4305] = 32'h248a57a2;
    ram_cell[    4306] = 32'h2d577c3c;
    ram_cell[    4307] = 32'h6116536f;
    ram_cell[    4308] = 32'h2e76ffa3;
    ram_cell[    4309] = 32'hdda2696a;
    ram_cell[    4310] = 32'he26a9f77;
    ram_cell[    4311] = 32'h8b66b017;
    ram_cell[    4312] = 32'hb1e61379;
    ram_cell[    4313] = 32'hc2eb16b4;
    ram_cell[    4314] = 32'h675b06fc;
    ram_cell[    4315] = 32'hfe67d891;
    ram_cell[    4316] = 32'h0879a9a6;
    ram_cell[    4317] = 32'h0085cee3;
    ram_cell[    4318] = 32'h5c1f12ce;
    ram_cell[    4319] = 32'h84e738c9;
    ram_cell[    4320] = 32'h32b423d4;
    ram_cell[    4321] = 32'hcf083d15;
    ram_cell[    4322] = 32'h8ca3971f;
    ram_cell[    4323] = 32'h15481fab;
    ram_cell[    4324] = 32'h2e0b1c56;
    ram_cell[    4325] = 32'h1f9ecda9;
    ram_cell[    4326] = 32'hfde4c5b1;
    ram_cell[    4327] = 32'hd7f31aad;
    ram_cell[    4328] = 32'hfd015a03;
    ram_cell[    4329] = 32'h9f4dccdc;
    ram_cell[    4330] = 32'h972d9dc9;
    ram_cell[    4331] = 32'h03153939;
    ram_cell[    4332] = 32'hcce37438;
    ram_cell[    4333] = 32'h89327be6;
    ram_cell[    4334] = 32'h6b02bcb8;
    ram_cell[    4335] = 32'ha87227a5;
    ram_cell[    4336] = 32'h7ab9cfca;
    ram_cell[    4337] = 32'hbbcd6450;
    ram_cell[    4338] = 32'h144d5c9c;
    ram_cell[    4339] = 32'hde280b01;
    ram_cell[    4340] = 32'h812c2eec;
    ram_cell[    4341] = 32'hc91d64ba;
    ram_cell[    4342] = 32'h5d717e00;
    ram_cell[    4343] = 32'hf0391f85;
    ram_cell[    4344] = 32'ha3cc5789;
    ram_cell[    4345] = 32'hd598ae7b;
    ram_cell[    4346] = 32'h7f4c6b2f;
    ram_cell[    4347] = 32'hc12abc39;
    ram_cell[    4348] = 32'haa58ee17;
    ram_cell[    4349] = 32'h90edeb07;
    ram_cell[    4350] = 32'h2b1e78c8;
    ram_cell[    4351] = 32'hed339580;
    ram_cell[    4352] = 32'h777d9b9a;
    ram_cell[    4353] = 32'h83402c7d;
    ram_cell[    4354] = 32'h7adfd76d;
    ram_cell[    4355] = 32'hf5bd1dac;
    ram_cell[    4356] = 32'hcaf73d13;
    ram_cell[    4357] = 32'h466f4e28;
    ram_cell[    4358] = 32'h8605d628;
    ram_cell[    4359] = 32'hd50d13cb;
    ram_cell[    4360] = 32'h99aa4e6b;
    ram_cell[    4361] = 32'h24a9083b;
    ram_cell[    4362] = 32'ha76aba58;
    ram_cell[    4363] = 32'he149be6c;
    ram_cell[    4364] = 32'h65db693d;
    ram_cell[    4365] = 32'h40aad0e1;
    ram_cell[    4366] = 32'h4b69c3ee;
    ram_cell[    4367] = 32'h757982a9;
    ram_cell[    4368] = 32'ha3cd6322;
    ram_cell[    4369] = 32'hb85e6d6f;
    ram_cell[    4370] = 32'hdba2a172;
    ram_cell[    4371] = 32'h45b50448;
    ram_cell[    4372] = 32'h255c599b;
    ram_cell[    4373] = 32'h8963ccd7;
    ram_cell[    4374] = 32'h9c7ef3ec;
    ram_cell[    4375] = 32'hf546c3fe;
    ram_cell[    4376] = 32'hcdc42853;
    ram_cell[    4377] = 32'h996c0c29;
    ram_cell[    4378] = 32'ha66a04a5;
    ram_cell[    4379] = 32'ha9909dea;
    ram_cell[    4380] = 32'hb517217a;
    ram_cell[    4381] = 32'h89dc536c;
    ram_cell[    4382] = 32'h25d73594;
    ram_cell[    4383] = 32'h891e67c2;
    ram_cell[    4384] = 32'h576c9b78;
    ram_cell[    4385] = 32'haac9899c;
    ram_cell[    4386] = 32'hab757489;
    ram_cell[    4387] = 32'h467be70c;
    ram_cell[    4388] = 32'h7bee1af6;
    ram_cell[    4389] = 32'h20e44198;
    ram_cell[    4390] = 32'h6c1b6513;
    ram_cell[    4391] = 32'hd491201e;
    ram_cell[    4392] = 32'hc0cd2896;
    ram_cell[    4393] = 32'hbbdcb179;
    ram_cell[    4394] = 32'h39b252df;
    ram_cell[    4395] = 32'h80863a0b;
    ram_cell[    4396] = 32'hdcf1974d;
    ram_cell[    4397] = 32'h72581231;
    ram_cell[    4398] = 32'ha56429e1;
    ram_cell[    4399] = 32'h80ff2218;
    ram_cell[    4400] = 32'hc3082207;
    ram_cell[    4401] = 32'h21ce05f9;
    ram_cell[    4402] = 32'hf21a7bdc;
    ram_cell[    4403] = 32'h48a1dff0;
    ram_cell[    4404] = 32'h5a774dc6;
    ram_cell[    4405] = 32'h04a54661;
    ram_cell[    4406] = 32'h63895d8b;
    ram_cell[    4407] = 32'h33e91d0f;
    ram_cell[    4408] = 32'h6a5a81a1;
    ram_cell[    4409] = 32'h853913fb;
    ram_cell[    4410] = 32'hc191c61a;
    ram_cell[    4411] = 32'h82d47a1d;
    ram_cell[    4412] = 32'hf442dc1d;
    ram_cell[    4413] = 32'h2d78b338;
    ram_cell[    4414] = 32'h5c48cf17;
    ram_cell[    4415] = 32'h95b9dcf5;
    ram_cell[    4416] = 32'h5d0d5960;
    ram_cell[    4417] = 32'h0f35dc36;
    ram_cell[    4418] = 32'h5d17722b;
    ram_cell[    4419] = 32'h3f0a01b4;
    ram_cell[    4420] = 32'h97c8ae34;
    ram_cell[    4421] = 32'h7e54eaeb;
    ram_cell[    4422] = 32'h31527db7;
    ram_cell[    4423] = 32'hda560ea4;
    ram_cell[    4424] = 32'h14eeebca;
    ram_cell[    4425] = 32'h8a4ab1dd;
    ram_cell[    4426] = 32'hc1677b7b;
    ram_cell[    4427] = 32'h25426931;
    ram_cell[    4428] = 32'h4b8cc9c0;
    ram_cell[    4429] = 32'h31a4bbac;
    ram_cell[    4430] = 32'h53c8392e;
    ram_cell[    4431] = 32'h7958ddd1;
    ram_cell[    4432] = 32'h6052bf27;
    ram_cell[    4433] = 32'hb46d5614;
    ram_cell[    4434] = 32'hcaa6b35a;
    ram_cell[    4435] = 32'hef626054;
    ram_cell[    4436] = 32'h2fa1c12c;
    ram_cell[    4437] = 32'h49ecf0dc;
    ram_cell[    4438] = 32'h1084172e;
    ram_cell[    4439] = 32'h8d7b18ee;
    ram_cell[    4440] = 32'h43f277cb;
    ram_cell[    4441] = 32'hc0b925d1;
    ram_cell[    4442] = 32'hb0bc8a24;
    ram_cell[    4443] = 32'h0e849704;
    ram_cell[    4444] = 32'h653c94c8;
    ram_cell[    4445] = 32'h69698c7d;
    ram_cell[    4446] = 32'h0da4b31f;
    ram_cell[    4447] = 32'hf4a7e6b1;
    ram_cell[    4448] = 32'hfa23c893;
    ram_cell[    4449] = 32'hdd49bb76;
    ram_cell[    4450] = 32'hadf57fbe;
    ram_cell[    4451] = 32'h85013649;
    ram_cell[    4452] = 32'h7f866e4f;
    ram_cell[    4453] = 32'h5adc3dcf;
    ram_cell[    4454] = 32'hcca4cfa8;
    ram_cell[    4455] = 32'h0e5afcc6;
    ram_cell[    4456] = 32'h5c153d82;
    ram_cell[    4457] = 32'h9398852d;
    ram_cell[    4458] = 32'hbbdd33fa;
    ram_cell[    4459] = 32'hfd558c25;
    ram_cell[    4460] = 32'hcfdb1da9;
    ram_cell[    4461] = 32'hd7037671;
    ram_cell[    4462] = 32'hff8bddf9;
    ram_cell[    4463] = 32'h60fdc966;
    ram_cell[    4464] = 32'h7c0e9b59;
    ram_cell[    4465] = 32'h51b053b0;
    ram_cell[    4466] = 32'hefaf0b8f;
    ram_cell[    4467] = 32'hf3801c37;
    ram_cell[    4468] = 32'hbdb1bde5;
    ram_cell[    4469] = 32'h5956d193;
    ram_cell[    4470] = 32'h8eb28911;
    ram_cell[    4471] = 32'h608b1858;
    ram_cell[    4472] = 32'he5a76ff8;
    ram_cell[    4473] = 32'hcd9c20e1;
    ram_cell[    4474] = 32'h87d7620e;
    ram_cell[    4475] = 32'hb745ca4b;
    ram_cell[    4476] = 32'h654fdc97;
    ram_cell[    4477] = 32'heab1e021;
    ram_cell[    4478] = 32'hd004c54d;
    ram_cell[    4479] = 32'hcadf5a55;
    ram_cell[    4480] = 32'hde5665b2;
    ram_cell[    4481] = 32'h33e1bc6c;
    ram_cell[    4482] = 32'h72f461a0;
    ram_cell[    4483] = 32'h0120f6b6;
    ram_cell[    4484] = 32'h15feab29;
    ram_cell[    4485] = 32'hcbc09776;
    ram_cell[    4486] = 32'hc6621e6a;
    ram_cell[    4487] = 32'h6f5f4ddc;
    ram_cell[    4488] = 32'h6be92274;
    ram_cell[    4489] = 32'h10a310d4;
    ram_cell[    4490] = 32'hc182e28a;
    ram_cell[    4491] = 32'hf1f01877;
    ram_cell[    4492] = 32'h0db862da;
    ram_cell[    4493] = 32'hfffeedf2;
    ram_cell[    4494] = 32'h56c0fb3d;
    ram_cell[    4495] = 32'h918cc421;
    ram_cell[    4496] = 32'h8ed9e26f;
    ram_cell[    4497] = 32'h98965f5e;
    ram_cell[    4498] = 32'he16df0bb;
    ram_cell[    4499] = 32'heb194960;
    ram_cell[    4500] = 32'he8d8dc65;
    ram_cell[    4501] = 32'h4832490a;
    ram_cell[    4502] = 32'hab3176e8;
    ram_cell[    4503] = 32'hc4949e83;
    ram_cell[    4504] = 32'h94e908f0;
    ram_cell[    4505] = 32'h5383ef29;
    ram_cell[    4506] = 32'h33f51609;
    ram_cell[    4507] = 32'hc7308496;
    ram_cell[    4508] = 32'h5361550c;
    ram_cell[    4509] = 32'h385c9ec7;
    ram_cell[    4510] = 32'h0e278516;
    ram_cell[    4511] = 32'h39f5d67a;
    ram_cell[    4512] = 32'hdc557f9c;
    ram_cell[    4513] = 32'hd32a4a4d;
    ram_cell[    4514] = 32'he9939871;
    ram_cell[    4515] = 32'hfeec2d78;
    ram_cell[    4516] = 32'hc0b44c79;
    ram_cell[    4517] = 32'h2b4d622b;
    ram_cell[    4518] = 32'h3c17d932;
    ram_cell[    4519] = 32'h7e17eb25;
    ram_cell[    4520] = 32'h6d08451e;
    ram_cell[    4521] = 32'h49db02ae;
    ram_cell[    4522] = 32'h41e42b19;
    ram_cell[    4523] = 32'h86fefefa;
    ram_cell[    4524] = 32'h84e08e1f;
    ram_cell[    4525] = 32'hfaf0129f;
    ram_cell[    4526] = 32'hca844ecc;
    ram_cell[    4527] = 32'h98bcda28;
    ram_cell[    4528] = 32'hac7e1504;
    ram_cell[    4529] = 32'hbda84038;
    ram_cell[    4530] = 32'h1fcce7a0;
    ram_cell[    4531] = 32'hb68ecc9a;
    ram_cell[    4532] = 32'h98a82119;
    ram_cell[    4533] = 32'h0f57df6b;
    ram_cell[    4534] = 32'h126d39e3;
    ram_cell[    4535] = 32'h8e48be6b;
    ram_cell[    4536] = 32'hb9679251;
    ram_cell[    4537] = 32'hcb1efed1;
    ram_cell[    4538] = 32'hdaee88be;
    ram_cell[    4539] = 32'h787ed0ca;
    ram_cell[    4540] = 32'h46a74128;
    ram_cell[    4541] = 32'h16bc45af;
    ram_cell[    4542] = 32'h3d8efec8;
    ram_cell[    4543] = 32'h13850403;
    ram_cell[    4544] = 32'h31340168;
    ram_cell[    4545] = 32'h0920d4c9;
    ram_cell[    4546] = 32'hef8e85c5;
    ram_cell[    4547] = 32'h29076c1b;
    ram_cell[    4548] = 32'h9dc05fe4;
    ram_cell[    4549] = 32'hd8d33c3a;
    ram_cell[    4550] = 32'hb1d37180;
    ram_cell[    4551] = 32'hbd263133;
    ram_cell[    4552] = 32'hb7f3c7d0;
    ram_cell[    4553] = 32'h78e89667;
    ram_cell[    4554] = 32'hb117c345;
    ram_cell[    4555] = 32'he8fd7dc9;
    ram_cell[    4556] = 32'h4643a11e;
    ram_cell[    4557] = 32'hce7f5ead;
    ram_cell[    4558] = 32'h6da69bfc;
    ram_cell[    4559] = 32'h066bd967;
    ram_cell[    4560] = 32'h625fc3a9;
    ram_cell[    4561] = 32'hb5201777;
    ram_cell[    4562] = 32'h0a59662d;
    ram_cell[    4563] = 32'h5febefeb;
    ram_cell[    4564] = 32'hcb265a7a;
    ram_cell[    4565] = 32'hb26daa9f;
    ram_cell[    4566] = 32'hfe84be8f;
    ram_cell[    4567] = 32'he78b45b2;
    ram_cell[    4568] = 32'h8d158f34;
    ram_cell[    4569] = 32'h85e50f4c;
    ram_cell[    4570] = 32'hf7d05208;
    ram_cell[    4571] = 32'h941c56a5;
    ram_cell[    4572] = 32'h1a6bd131;
    ram_cell[    4573] = 32'h954255b0;
    ram_cell[    4574] = 32'h9a2703b5;
    ram_cell[    4575] = 32'h86dd809d;
    ram_cell[    4576] = 32'h1b8c6838;
    ram_cell[    4577] = 32'h6e36859c;
    ram_cell[    4578] = 32'h9189f233;
    ram_cell[    4579] = 32'h1c52e8b6;
    ram_cell[    4580] = 32'h3abff25e;
    ram_cell[    4581] = 32'h49de0a6c;
    ram_cell[    4582] = 32'h18ec3b15;
    ram_cell[    4583] = 32'h4bbf0d6b;
    ram_cell[    4584] = 32'h15dfbc3a;
    ram_cell[    4585] = 32'h380c267c;
    ram_cell[    4586] = 32'h004bab95;
    ram_cell[    4587] = 32'h34c0628f;
    ram_cell[    4588] = 32'h244b69d4;
    ram_cell[    4589] = 32'h9dec79ab;
    ram_cell[    4590] = 32'ha38b5e05;
    ram_cell[    4591] = 32'h630046de;
    ram_cell[    4592] = 32'ha618e99a;
    ram_cell[    4593] = 32'h88ece3d0;
    ram_cell[    4594] = 32'h1ce66e98;
    ram_cell[    4595] = 32'h746f1e30;
    ram_cell[    4596] = 32'h23a53fb9;
    ram_cell[    4597] = 32'hcc2ae09b;
    ram_cell[    4598] = 32'hf997cfc4;
    ram_cell[    4599] = 32'hbb9361c9;
    ram_cell[    4600] = 32'hd734bf5f;
    ram_cell[    4601] = 32'hbc86cc5d;
    ram_cell[    4602] = 32'h9fc5c0c9;
    ram_cell[    4603] = 32'h6189ac46;
    ram_cell[    4604] = 32'h0e2d4c90;
    ram_cell[    4605] = 32'h0fcba036;
    ram_cell[    4606] = 32'h58996c85;
    ram_cell[    4607] = 32'h5d20b768;
    ram_cell[    4608] = 32'heb9a4c92;
    ram_cell[    4609] = 32'h1be69113;
    ram_cell[    4610] = 32'h7ca0a7a3;
    ram_cell[    4611] = 32'h96fa9a10;
    ram_cell[    4612] = 32'h1cbce2b1;
    ram_cell[    4613] = 32'hc55f4ddd;
    ram_cell[    4614] = 32'h84caaa94;
    ram_cell[    4615] = 32'h4f068af8;
    ram_cell[    4616] = 32'h622d154b;
    ram_cell[    4617] = 32'hd40e346e;
    ram_cell[    4618] = 32'h3af6c50f;
    ram_cell[    4619] = 32'h5a50c821;
    ram_cell[    4620] = 32'h43f9620f;
    ram_cell[    4621] = 32'h32e05534;
    ram_cell[    4622] = 32'h94613066;
    ram_cell[    4623] = 32'h47f611a7;
    ram_cell[    4624] = 32'h94495510;
    ram_cell[    4625] = 32'h69af0eb8;
    ram_cell[    4626] = 32'h9f3eec43;
    ram_cell[    4627] = 32'h7ba65d4b;
    ram_cell[    4628] = 32'h2999cac8;
    ram_cell[    4629] = 32'h2b56ded1;
    ram_cell[    4630] = 32'hfa0fe5fd;
    ram_cell[    4631] = 32'h6e54858f;
    ram_cell[    4632] = 32'h24246682;
    ram_cell[    4633] = 32'he0dbe528;
    ram_cell[    4634] = 32'ha441fa9a;
    ram_cell[    4635] = 32'ha82b65a9;
    ram_cell[    4636] = 32'ha1256b28;
    ram_cell[    4637] = 32'ha15d1e0c;
    ram_cell[    4638] = 32'h0e57036e;
    ram_cell[    4639] = 32'h60b65d37;
    ram_cell[    4640] = 32'hfa0dbf88;
    ram_cell[    4641] = 32'hc918479d;
    ram_cell[    4642] = 32'h49f80e47;
    ram_cell[    4643] = 32'h47255525;
    ram_cell[    4644] = 32'h2220d74c;
    ram_cell[    4645] = 32'h4ac411ef;
    ram_cell[    4646] = 32'h1a8935f9;
    ram_cell[    4647] = 32'h542abdcd;
    ram_cell[    4648] = 32'h85845969;
    ram_cell[    4649] = 32'hbb61d75f;
    ram_cell[    4650] = 32'hb951a2f9;
    ram_cell[    4651] = 32'h66c0cb8b;
    ram_cell[    4652] = 32'h9548cb64;
    ram_cell[    4653] = 32'ha99758a5;
    ram_cell[    4654] = 32'hb49f6106;
    ram_cell[    4655] = 32'h97c2d796;
    ram_cell[    4656] = 32'h691d8b3c;
    ram_cell[    4657] = 32'h71cdf105;
    ram_cell[    4658] = 32'h4897eb84;
    ram_cell[    4659] = 32'h58a4a0ac;
    ram_cell[    4660] = 32'hdc70cb20;
    ram_cell[    4661] = 32'h898f0ff4;
    ram_cell[    4662] = 32'h36ee86f9;
    ram_cell[    4663] = 32'h14198fec;
    ram_cell[    4664] = 32'h18c65a8b;
    ram_cell[    4665] = 32'hb6ba4601;
    ram_cell[    4666] = 32'h5e3f32f9;
    ram_cell[    4667] = 32'h098319ca;
    ram_cell[    4668] = 32'h0a23cd1d;
    ram_cell[    4669] = 32'h43654028;
    ram_cell[    4670] = 32'h1cbc66f5;
    ram_cell[    4671] = 32'hb7bd9e50;
    ram_cell[    4672] = 32'h73611c06;
    ram_cell[    4673] = 32'h48370fa6;
    ram_cell[    4674] = 32'hdc932f99;
    ram_cell[    4675] = 32'h1651a85a;
    ram_cell[    4676] = 32'hcd7c0916;
    ram_cell[    4677] = 32'h946cfa99;
    ram_cell[    4678] = 32'h82a7b1cd;
    ram_cell[    4679] = 32'ha0e866ed;
    ram_cell[    4680] = 32'h95e2e99e;
    ram_cell[    4681] = 32'he999144c;
    ram_cell[    4682] = 32'h1e78acf5;
    ram_cell[    4683] = 32'h63dc5714;
    ram_cell[    4684] = 32'hf59975d6;
    ram_cell[    4685] = 32'h15826c61;
    ram_cell[    4686] = 32'he5ed8720;
    ram_cell[    4687] = 32'h1645a0cc;
    ram_cell[    4688] = 32'hd0b151eb;
    ram_cell[    4689] = 32'hbfc99e69;
    ram_cell[    4690] = 32'hc063f4cc;
    ram_cell[    4691] = 32'h52c5bf3e;
    ram_cell[    4692] = 32'hccb1d2fd;
    ram_cell[    4693] = 32'h08a77229;
    ram_cell[    4694] = 32'he366361e;
    ram_cell[    4695] = 32'h810544a4;
    ram_cell[    4696] = 32'h3319cf86;
    ram_cell[    4697] = 32'h2e128a7a;
    ram_cell[    4698] = 32'hd42a24ca;
    ram_cell[    4699] = 32'hac2ca88e;
    ram_cell[    4700] = 32'hf8305576;
    ram_cell[    4701] = 32'h86088a74;
    ram_cell[    4702] = 32'h3a28c3ee;
    ram_cell[    4703] = 32'h5c8f77bf;
    ram_cell[    4704] = 32'h0447410c;
    ram_cell[    4705] = 32'h039af7b5;
    ram_cell[    4706] = 32'h6624ac85;
    ram_cell[    4707] = 32'hc505c630;
    ram_cell[    4708] = 32'h0a693910;
    ram_cell[    4709] = 32'hb95a52d2;
    ram_cell[    4710] = 32'h1ce56083;
    ram_cell[    4711] = 32'h3bddc2a7;
    ram_cell[    4712] = 32'h14e1dd96;
    ram_cell[    4713] = 32'he8569a0b;
    ram_cell[    4714] = 32'h6ff6ac85;
    ram_cell[    4715] = 32'hd94bd3d1;
    ram_cell[    4716] = 32'h8781db5c;
    ram_cell[    4717] = 32'h526ce9e2;
    ram_cell[    4718] = 32'hd1bef95e;
    ram_cell[    4719] = 32'h7c6b4be2;
    ram_cell[    4720] = 32'he31f81a1;
    ram_cell[    4721] = 32'h553e5f09;
    ram_cell[    4722] = 32'h973c6a1a;
    ram_cell[    4723] = 32'h31333818;
    ram_cell[    4724] = 32'h7ef00708;
    ram_cell[    4725] = 32'h6033213b;
    ram_cell[    4726] = 32'h4edcd83a;
    ram_cell[    4727] = 32'h31f5e049;
    ram_cell[    4728] = 32'h17f50a05;
    ram_cell[    4729] = 32'h84b0ed58;
    ram_cell[    4730] = 32'hb5fc335b;
    ram_cell[    4731] = 32'h297c6dd3;
    ram_cell[    4732] = 32'hb7e2c805;
    ram_cell[    4733] = 32'h8f6c12af;
    ram_cell[    4734] = 32'h4ce848c2;
    ram_cell[    4735] = 32'h746a6218;
    ram_cell[    4736] = 32'h90d8e540;
    ram_cell[    4737] = 32'h705c5691;
    ram_cell[    4738] = 32'hd7004684;
    ram_cell[    4739] = 32'h3026c3a3;
    ram_cell[    4740] = 32'h6cfe702e;
    ram_cell[    4741] = 32'h5955c62a;
    ram_cell[    4742] = 32'hf266add2;
    ram_cell[    4743] = 32'h7cb4c3d8;
    ram_cell[    4744] = 32'h7e18b23e;
    ram_cell[    4745] = 32'h7ac1bf90;
    ram_cell[    4746] = 32'he0e25978;
    ram_cell[    4747] = 32'h7035627a;
    ram_cell[    4748] = 32'hfab8ce5b;
    ram_cell[    4749] = 32'ha1cf3844;
    ram_cell[    4750] = 32'h88382442;
    ram_cell[    4751] = 32'h95f7bdcd;
    ram_cell[    4752] = 32'he1534bce;
    ram_cell[    4753] = 32'hd5cdf400;
    ram_cell[    4754] = 32'h240aacc0;
    ram_cell[    4755] = 32'h3e9d612d;
    ram_cell[    4756] = 32'h9e2c1a8a;
    ram_cell[    4757] = 32'h6995bf65;
    ram_cell[    4758] = 32'h560f0632;
    ram_cell[    4759] = 32'hf7a72b8e;
    ram_cell[    4760] = 32'he091eb92;
    ram_cell[    4761] = 32'hf02c2c74;
    ram_cell[    4762] = 32'h8096cb04;
    ram_cell[    4763] = 32'h6457b082;
    ram_cell[    4764] = 32'h777477cc;
    ram_cell[    4765] = 32'h4e7ffc16;
    ram_cell[    4766] = 32'haabfe5de;
    ram_cell[    4767] = 32'hc189520b;
    ram_cell[    4768] = 32'h31e80bf2;
    ram_cell[    4769] = 32'h46905134;
    ram_cell[    4770] = 32'h5293feba;
    ram_cell[    4771] = 32'h3998abc6;
    ram_cell[    4772] = 32'h780ce118;
    ram_cell[    4773] = 32'hfe83a5d8;
    ram_cell[    4774] = 32'h773088f0;
    ram_cell[    4775] = 32'hff92be7d;
    ram_cell[    4776] = 32'h04eead46;
    ram_cell[    4777] = 32'h1213462c;
    ram_cell[    4778] = 32'h72ff5caf;
    ram_cell[    4779] = 32'hd55f089d;
    ram_cell[    4780] = 32'h8654d412;
    ram_cell[    4781] = 32'hb31734ee;
    ram_cell[    4782] = 32'h9f94935e;
    ram_cell[    4783] = 32'h69e1ebb3;
    ram_cell[    4784] = 32'he381715a;
    ram_cell[    4785] = 32'h8a53ff38;
    ram_cell[    4786] = 32'h9431c527;
    ram_cell[    4787] = 32'h1510cc73;
    ram_cell[    4788] = 32'h538c3493;
    ram_cell[    4789] = 32'h46f750df;
    ram_cell[    4790] = 32'hb3db3f98;
    ram_cell[    4791] = 32'ha0453af5;
    ram_cell[    4792] = 32'h0d8f8617;
    ram_cell[    4793] = 32'h8f31ba9e;
    ram_cell[    4794] = 32'hc5a1ce89;
    ram_cell[    4795] = 32'hdde371e3;
    ram_cell[    4796] = 32'h34b855de;
    ram_cell[    4797] = 32'hf87cdb35;
    ram_cell[    4798] = 32'hc502a164;
    ram_cell[    4799] = 32'h9b6ffefd;
    ram_cell[    4800] = 32'hac16923c;
    ram_cell[    4801] = 32'h85855421;
    ram_cell[    4802] = 32'h67f64600;
    ram_cell[    4803] = 32'h040e08da;
    ram_cell[    4804] = 32'h22b406fa;
    ram_cell[    4805] = 32'h38850cc4;
    ram_cell[    4806] = 32'h33a6bd67;
    ram_cell[    4807] = 32'h64b6304b;
    ram_cell[    4808] = 32'hdd94005f;
    ram_cell[    4809] = 32'hcd195842;
    ram_cell[    4810] = 32'h5f1abc79;
    ram_cell[    4811] = 32'h188ff238;
    ram_cell[    4812] = 32'h1930838a;
    ram_cell[    4813] = 32'h95eb904a;
    ram_cell[    4814] = 32'hcb366872;
    ram_cell[    4815] = 32'hba970b41;
    ram_cell[    4816] = 32'h73dd9d96;
    ram_cell[    4817] = 32'h31fc0dfd;
    ram_cell[    4818] = 32'h6ab0f6bf;
    ram_cell[    4819] = 32'h33d0873e;
    ram_cell[    4820] = 32'h1dcfc9c4;
    ram_cell[    4821] = 32'h8b279192;
    ram_cell[    4822] = 32'h441a29d6;
    ram_cell[    4823] = 32'h07777f99;
    ram_cell[    4824] = 32'h5b4ccb28;
    ram_cell[    4825] = 32'h231f0d2e;
    ram_cell[    4826] = 32'h7003b804;
    ram_cell[    4827] = 32'hf882c398;
    ram_cell[    4828] = 32'h0fbb2c30;
    ram_cell[    4829] = 32'h14ad591b;
    ram_cell[    4830] = 32'hdbede1c2;
    ram_cell[    4831] = 32'hea74007d;
    ram_cell[    4832] = 32'h5bbd0186;
    ram_cell[    4833] = 32'hb5c18b1a;
    ram_cell[    4834] = 32'h865e45de;
    ram_cell[    4835] = 32'h209ceb67;
    ram_cell[    4836] = 32'h31edd65a;
    ram_cell[    4837] = 32'h779fec11;
    ram_cell[    4838] = 32'h02235599;
    ram_cell[    4839] = 32'hfcb46719;
    ram_cell[    4840] = 32'hfb8b9520;
    ram_cell[    4841] = 32'hcdbe5f51;
    ram_cell[    4842] = 32'h41772178;
    ram_cell[    4843] = 32'h5676d8b7;
    ram_cell[    4844] = 32'h83f2a470;
    ram_cell[    4845] = 32'h3a11d7ed;
    ram_cell[    4846] = 32'hc7b892cf;
    ram_cell[    4847] = 32'h8c80199d;
    ram_cell[    4848] = 32'h80460e05;
    ram_cell[    4849] = 32'h0d8095a4;
    ram_cell[    4850] = 32'h8687b768;
    ram_cell[    4851] = 32'ha5795b9f;
    ram_cell[    4852] = 32'h38d0d2bf;
    ram_cell[    4853] = 32'hb0db1d2c;
    ram_cell[    4854] = 32'he6dbb953;
    ram_cell[    4855] = 32'h1a0111bd;
    ram_cell[    4856] = 32'h25ca4e91;
    ram_cell[    4857] = 32'h372816d6;
    ram_cell[    4858] = 32'h5012cf10;
    ram_cell[    4859] = 32'h891a22f8;
    ram_cell[    4860] = 32'hc8e460ef;
    ram_cell[    4861] = 32'h2ce93eed;
    ram_cell[    4862] = 32'h400730bc;
    ram_cell[    4863] = 32'h597c58c8;
    ram_cell[    4864] = 32'hd3254c20;
    ram_cell[    4865] = 32'h425accc2;
    ram_cell[    4866] = 32'h1ae52af1;
    ram_cell[    4867] = 32'hd829ce61;
    ram_cell[    4868] = 32'h8f211065;
    ram_cell[    4869] = 32'hc53976c5;
    ram_cell[    4870] = 32'hf0781d46;
    ram_cell[    4871] = 32'hbe14a4a7;
    ram_cell[    4872] = 32'hbe83750b;
    ram_cell[    4873] = 32'h57c540e6;
    ram_cell[    4874] = 32'h51ba9d4e;
    ram_cell[    4875] = 32'hca74d7e8;
    ram_cell[    4876] = 32'h00844220;
    ram_cell[    4877] = 32'he6d09304;
    ram_cell[    4878] = 32'h0d2aa452;
    ram_cell[    4879] = 32'hd6e986f4;
    ram_cell[    4880] = 32'h70dc1238;
    ram_cell[    4881] = 32'h143b6b0e;
    ram_cell[    4882] = 32'h23206817;
    ram_cell[    4883] = 32'h826348c8;
    ram_cell[    4884] = 32'hd5f9a82c;
    ram_cell[    4885] = 32'h4c746134;
    ram_cell[    4886] = 32'h09a27b19;
    ram_cell[    4887] = 32'h03fb36fe;
    ram_cell[    4888] = 32'h1655c9b9;
    ram_cell[    4889] = 32'h31e9b4a4;
    ram_cell[    4890] = 32'h6f1ccf61;
    ram_cell[    4891] = 32'h1271f07a;
    ram_cell[    4892] = 32'hc3779640;
    ram_cell[    4893] = 32'hb20e17e7;
    ram_cell[    4894] = 32'h01f54e60;
    ram_cell[    4895] = 32'h8c3f8398;
    ram_cell[    4896] = 32'hfd1a3966;
    ram_cell[    4897] = 32'h26994dd8;
    ram_cell[    4898] = 32'hd0811d40;
    ram_cell[    4899] = 32'hdb5d399c;
    ram_cell[    4900] = 32'h40970242;
    ram_cell[    4901] = 32'hf6fca543;
    ram_cell[    4902] = 32'h836bdaa7;
    ram_cell[    4903] = 32'h97457044;
    ram_cell[    4904] = 32'hcaf8e8cc;
    ram_cell[    4905] = 32'h201afc25;
    ram_cell[    4906] = 32'hfd8ec878;
    ram_cell[    4907] = 32'he55c2e1b;
    ram_cell[    4908] = 32'hb29d4c37;
    ram_cell[    4909] = 32'h88b106a9;
    ram_cell[    4910] = 32'h168f8c22;
    ram_cell[    4911] = 32'hc2401b53;
    ram_cell[    4912] = 32'h74186e75;
    ram_cell[    4913] = 32'h8468e87a;
    ram_cell[    4914] = 32'hb4b2a101;
    ram_cell[    4915] = 32'hfe7367a2;
    ram_cell[    4916] = 32'h808b5dc1;
    ram_cell[    4917] = 32'h764caa46;
    ram_cell[    4918] = 32'hf29590c2;
    ram_cell[    4919] = 32'h81e32ffb;
    ram_cell[    4920] = 32'h28358cc2;
    ram_cell[    4921] = 32'h099396ec;
    ram_cell[    4922] = 32'h009553e7;
    ram_cell[    4923] = 32'h2764b3b0;
    ram_cell[    4924] = 32'he4fee560;
    ram_cell[    4925] = 32'h4e7cd1a6;
    ram_cell[    4926] = 32'h039794a8;
    ram_cell[    4927] = 32'hbf0f75cb;
    ram_cell[    4928] = 32'h39e0fb3b;
    ram_cell[    4929] = 32'h559361ed;
    ram_cell[    4930] = 32'hcffdcc12;
    ram_cell[    4931] = 32'h4e6ae2a2;
    ram_cell[    4932] = 32'hd702a841;
    ram_cell[    4933] = 32'h2d3467d9;
    ram_cell[    4934] = 32'hc2000a7c;
    ram_cell[    4935] = 32'h057875ec;
    ram_cell[    4936] = 32'h9d08e52c;
    ram_cell[    4937] = 32'h48445861;
    ram_cell[    4938] = 32'h6001d008;
    ram_cell[    4939] = 32'hf3a92a09;
    ram_cell[    4940] = 32'h751f9065;
    ram_cell[    4941] = 32'h900c8d32;
    ram_cell[    4942] = 32'hd6e27357;
    ram_cell[    4943] = 32'hc2f10eb7;
    ram_cell[    4944] = 32'hc1c2ff1d;
    ram_cell[    4945] = 32'h04b10353;
    ram_cell[    4946] = 32'h32d17687;
    ram_cell[    4947] = 32'h07c667ce;
    ram_cell[    4948] = 32'hb7b80989;
    ram_cell[    4949] = 32'h0db6a739;
    ram_cell[    4950] = 32'h2c7a4cdd;
    ram_cell[    4951] = 32'hafcf5401;
    ram_cell[    4952] = 32'hfe82c50b;
    ram_cell[    4953] = 32'h05d649a7;
    ram_cell[    4954] = 32'he97d693d;
    ram_cell[    4955] = 32'he109ef0d;
    ram_cell[    4956] = 32'hd5ad8b35;
    ram_cell[    4957] = 32'h579b93bb;
    ram_cell[    4958] = 32'h66ceaf45;
    ram_cell[    4959] = 32'h8368fa4f;
    ram_cell[    4960] = 32'hdf27f990;
    ram_cell[    4961] = 32'hba7d3d92;
    ram_cell[    4962] = 32'hb24546de;
    ram_cell[    4963] = 32'h1b73a4e2;
    ram_cell[    4964] = 32'ha6dbda15;
    ram_cell[    4965] = 32'hcb120d31;
    ram_cell[    4966] = 32'hc47a8723;
    ram_cell[    4967] = 32'hd6930447;
    ram_cell[    4968] = 32'haf1606d7;
    ram_cell[    4969] = 32'h80c122ea;
    ram_cell[    4970] = 32'h3f7cefaa;
    ram_cell[    4971] = 32'h8ff5a481;
    ram_cell[    4972] = 32'h0801eb47;
    ram_cell[    4973] = 32'h7c4a13ec;
    ram_cell[    4974] = 32'h4c9017fa;
    ram_cell[    4975] = 32'hbaeacaa6;
    ram_cell[    4976] = 32'ha1c46cda;
    ram_cell[    4977] = 32'h3f577c02;
    ram_cell[    4978] = 32'h8e35716a;
    ram_cell[    4979] = 32'h26e42306;
    ram_cell[    4980] = 32'h1fad32cc;
    ram_cell[    4981] = 32'h6c29ae09;
    ram_cell[    4982] = 32'h0392e831;
    ram_cell[    4983] = 32'h728d0e5e;
    ram_cell[    4984] = 32'hb6ac2cfa;
    ram_cell[    4985] = 32'h93b04bac;
    ram_cell[    4986] = 32'h7760c3d9;
    ram_cell[    4987] = 32'h53ec680f;
    ram_cell[    4988] = 32'h915af0de;
    ram_cell[    4989] = 32'hba844e2a;
    ram_cell[    4990] = 32'hec772c28;
    ram_cell[    4991] = 32'h42a61263;
    ram_cell[    4992] = 32'h0aa6aaec;
    ram_cell[    4993] = 32'h4186b296;
    ram_cell[    4994] = 32'h6d0618ce;
    ram_cell[    4995] = 32'h2c5c5539;
    ram_cell[    4996] = 32'h18233ab3;
    ram_cell[    4997] = 32'h69ee9053;
    ram_cell[    4998] = 32'h191a78a2;
    ram_cell[    4999] = 32'h2a0aa9bc;
    ram_cell[    5000] = 32'h3aabd964;
    ram_cell[    5001] = 32'hcc766326;
    ram_cell[    5002] = 32'hb3ef01cf;
    ram_cell[    5003] = 32'hfb89a5e8;
    ram_cell[    5004] = 32'hf0a75c01;
    ram_cell[    5005] = 32'hb6789423;
    ram_cell[    5006] = 32'h645470f5;
    ram_cell[    5007] = 32'hed60c64a;
    ram_cell[    5008] = 32'hdc27f56c;
    ram_cell[    5009] = 32'hdd0132a7;
    ram_cell[    5010] = 32'he9b21c06;
    ram_cell[    5011] = 32'hfcfe3310;
    ram_cell[    5012] = 32'hb480fb98;
    ram_cell[    5013] = 32'ha2131617;
    ram_cell[    5014] = 32'h11b9d61d;
    ram_cell[    5015] = 32'h592cebf3;
    ram_cell[    5016] = 32'h5f657cfb;
    ram_cell[    5017] = 32'h170a7589;
    ram_cell[    5018] = 32'ha0b899f3;
    ram_cell[    5019] = 32'h2dddfe78;
    ram_cell[    5020] = 32'h9ad8b08f;
    ram_cell[    5021] = 32'hd33a5836;
    ram_cell[    5022] = 32'ha7eb22d3;
    ram_cell[    5023] = 32'ha8c9cd5a;
    ram_cell[    5024] = 32'hb53e5de5;
    ram_cell[    5025] = 32'he03355e4;
    ram_cell[    5026] = 32'hd161e0c8;
    ram_cell[    5027] = 32'h35102b6d;
    ram_cell[    5028] = 32'h43acecff;
    ram_cell[    5029] = 32'hdbb634f7;
    ram_cell[    5030] = 32'h34930bdd;
    ram_cell[    5031] = 32'h695e796e;
    ram_cell[    5032] = 32'h4c7b457f;
    ram_cell[    5033] = 32'h69b7796e;
    ram_cell[    5034] = 32'h6ec1058d;
    ram_cell[    5035] = 32'h07ee4d8f;
    ram_cell[    5036] = 32'h22c8ca3e;
    ram_cell[    5037] = 32'h16cb9f4d;
    ram_cell[    5038] = 32'hf18a587b;
    ram_cell[    5039] = 32'h3eb1b952;
    ram_cell[    5040] = 32'h99b86b77;
    ram_cell[    5041] = 32'h13ab8041;
    ram_cell[    5042] = 32'hfe417445;
    ram_cell[    5043] = 32'h98848d77;
    ram_cell[    5044] = 32'he619bd79;
    ram_cell[    5045] = 32'h0ce0fe9b;
    ram_cell[    5046] = 32'h7eba2676;
    ram_cell[    5047] = 32'hb560287c;
    ram_cell[    5048] = 32'h2007282a;
    ram_cell[    5049] = 32'h09ee043b;
    ram_cell[    5050] = 32'h7aaa4542;
    ram_cell[    5051] = 32'ha00c271f;
    ram_cell[    5052] = 32'h8b466508;
    ram_cell[    5053] = 32'h19cfc188;
    ram_cell[    5054] = 32'h606a355d;
    ram_cell[    5055] = 32'h839e83c4;
    ram_cell[    5056] = 32'h9e6dc676;
    ram_cell[    5057] = 32'h4fde88e4;
    ram_cell[    5058] = 32'h0d976419;
    ram_cell[    5059] = 32'hfb2aaf0a;
    ram_cell[    5060] = 32'h5b2964e2;
    ram_cell[    5061] = 32'h0e6f010c;
    ram_cell[    5062] = 32'hc165fcee;
    ram_cell[    5063] = 32'h370d96d4;
    ram_cell[    5064] = 32'hf1f17926;
    ram_cell[    5065] = 32'h36d3f41a;
    ram_cell[    5066] = 32'hade739a0;
    ram_cell[    5067] = 32'h85556736;
    ram_cell[    5068] = 32'h561b735a;
    ram_cell[    5069] = 32'hdebb1172;
    ram_cell[    5070] = 32'h388fc43a;
    ram_cell[    5071] = 32'h82cee0c9;
    ram_cell[    5072] = 32'h9e402d0b;
    ram_cell[    5073] = 32'hfa056831;
    ram_cell[    5074] = 32'hdd3f04d3;
    ram_cell[    5075] = 32'h3b024467;
    ram_cell[    5076] = 32'h9e79fb77;
    ram_cell[    5077] = 32'h6ada23c7;
    ram_cell[    5078] = 32'hca786f6a;
    ram_cell[    5079] = 32'h63ef4a1a;
    ram_cell[    5080] = 32'hb8179cb8;
    ram_cell[    5081] = 32'hefa64b49;
    ram_cell[    5082] = 32'h60a9d6be;
    ram_cell[    5083] = 32'h64505926;
    ram_cell[    5084] = 32'hd109f3ad;
    ram_cell[    5085] = 32'hd5177071;
    ram_cell[    5086] = 32'hcc39e0e5;
    ram_cell[    5087] = 32'hef34ebbc;
    ram_cell[    5088] = 32'h7b865ba3;
    ram_cell[    5089] = 32'h5658a98a;
    ram_cell[    5090] = 32'hd198895a;
    ram_cell[    5091] = 32'h8b99106c;
    ram_cell[    5092] = 32'h919f9591;
    ram_cell[    5093] = 32'h68668e12;
    ram_cell[    5094] = 32'h41111576;
    ram_cell[    5095] = 32'h9d36048e;
    ram_cell[    5096] = 32'hed255768;
    ram_cell[    5097] = 32'h9f0352ee;
    ram_cell[    5098] = 32'hdc329f16;
    ram_cell[    5099] = 32'h5807d306;
    ram_cell[    5100] = 32'hb37fc7e4;
    ram_cell[    5101] = 32'h728b63af;
    ram_cell[    5102] = 32'h1c602528;
    ram_cell[    5103] = 32'h68c28349;
    ram_cell[    5104] = 32'hdb804b31;
    ram_cell[    5105] = 32'h5a1c665b;
    ram_cell[    5106] = 32'hfc8aa90c;
    ram_cell[    5107] = 32'hfce34008;
    ram_cell[    5108] = 32'h9c5e2951;
    ram_cell[    5109] = 32'hcb728f98;
    ram_cell[    5110] = 32'h80b1b97c;
    ram_cell[    5111] = 32'hd63932aa;
    ram_cell[    5112] = 32'hd772ada5;
    ram_cell[    5113] = 32'hd27b0d79;
    ram_cell[    5114] = 32'he48755a4;
    ram_cell[    5115] = 32'he8df21bf;
    ram_cell[    5116] = 32'he46b3fd4;
    ram_cell[    5117] = 32'h1b50669b;
    ram_cell[    5118] = 32'h443b893c;
    ram_cell[    5119] = 32'h92ff2c6f;
    ram_cell[    5120] = 32'hb7096856;
    ram_cell[    5121] = 32'h89510dbb;
    ram_cell[    5122] = 32'h7bbc61f2;
    ram_cell[    5123] = 32'hb108deca;
    ram_cell[    5124] = 32'h832c96a1;
    ram_cell[    5125] = 32'hd4c8de74;
    ram_cell[    5126] = 32'h33312733;
    ram_cell[    5127] = 32'ha952a460;
    ram_cell[    5128] = 32'h8f797b9c;
    ram_cell[    5129] = 32'h52dfa82a;
    ram_cell[    5130] = 32'hfd6dd371;
    ram_cell[    5131] = 32'h8a9b0045;
    ram_cell[    5132] = 32'hf2dfadf6;
    ram_cell[    5133] = 32'h4869a48d;
    ram_cell[    5134] = 32'h7f81309f;
    ram_cell[    5135] = 32'h7b6ec299;
    ram_cell[    5136] = 32'hce7bd6c9;
    ram_cell[    5137] = 32'hbb512bff;
    ram_cell[    5138] = 32'h7575d494;
    ram_cell[    5139] = 32'h693a60bd;
    ram_cell[    5140] = 32'hae371f5e;
    ram_cell[    5141] = 32'h4f1524a6;
    ram_cell[    5142] = 32'h29d933b6;
    ram_cell[    5143] = 32'heba15003;
    ram_cell[    5144] = 32'hb068e087;
    ram_cell[    5145] = 32'h656d4105;
    ram_cell[    5146] = 32'h9b499537;
    ram_cell[    5147] = 32'hbfc48a52;
    ram_cell[    5148] = 32'h0f86659b;
    ram_cell[    5149] = 32'hec83764b;
    ram_cell[    5150] = 32'h63b25108;
    ram_cell[    5151] = 32'hd99492b5;
    ram_cell[    5152] = 32'h61e7ad52;
    ram_cell[    5153] = 32'h0a44a547;
    ram_cell[    5154] = 32'h39d00cd7;
    ram_cell[    5155] = 32'h0cdfc7f6;
    ram_cell[    5156] = 32'h243e9011;
    ram_cell[    5157] = 32'h725a964d;
    ram_cell[    5158] = 32'h68ae2b12;
    ram_cell[    5159] = 32'hc9c11f9f;
    ram_cell[    5160] = 32'he28e4c43;
    ram_cell[    5161] = 32'hfb1f2885;
    ram_cell[    5162] = 32'hcba1f1f4;
    ram_cell[    5163] = 32'ha9f98930;
    ram_cell[    5164] = 32'h32ea0d65;
    ram_cell[    5165] = 32'h92b2f38a;
    ram_cell[    5166] = 32'h65511a18;
    ram_cell[    5167] = 32'hdb805551;
    ram_cell[    5168] = 32'h98791d2c;
    ram_cell[    5169] = 32'hc57289cd;
    ram_cell[    5170] = 32'hec250b35;
    ram_cell[    5171] = 32'hd7fa3fc7;
    ram_cell[    5172] = 32'hc642ae6c;
    ram_cell[    5173] = 32'h7e72e104;
    ram_cell[    5174] = 32'h50cc0098;
    ram_cell[    5175] = 32'h23d5cad7;
    ram_cell[    5176] = 32'h07839ca7;
    ram_cell[    5177] = 32'he3d5ad65;
    ram_cell[    5178] = 32'h5e4f3e1b;
    ram_cell[    5179] = 32'heff9646a;
    ram_cell[    5180] = 32'hf163c50d;
    ram_cell[    5181] = 32'h4a16e46b;
    ram_cell[    5182] = 32'h49504508;
    ram_cell[    5183] = 32'h6f2b1b41;
    ram_cell[    5184] = 32'h4566fc37;
    ram_cell[    5185] = 32'h5d812bc8;
    ram_cell[    5186] = 32'he569edc3;
    ram_cell[    5187] = 32'hac1ec6ed;
    ram_cell[    5188] = 32'h642f807e;
    ram_cell[    5189] = 32'hf2da1f63;
    ram_cell[    5190] = 32'h2640560a;
    ram_cell[    5191] = 32'ha30c535f;
    ram_cell[    5192] = 32'h82ba6ee3;
    ram_cell[    5193] = 32'h20c9be0a;
    ram_cell[    5194] = 32'hac4c7c72;
    ram_cell[    5195] = 32'hf31ab09c;
    ram_cell[    5196] = 32'h768979e6;
    ram_cell[    5197] = 32'h3694ff6b;
    ram_cell[    5198] = 32'habe5feda;
    ram_cell[    5199] = 32'h93399740;
    ram_cell[    5200] = 32'h490dffd2;
    ram_cell[    5201] = 32'hc8245128;
    ram_cell[    5202] = 32'h421f2ae3;
    ram_cell[    5203] = 32'h68be0f47;
    ram_cell[    5204] = 32'h0ba93d01;
    ram_cell[    5205] = 32'h1388c594;
    ram_cell[    5206] = 32'he8a62831;
    ram_cell[    5207] = 32'h20102570;
    ram_cell[    5208] = 32'h7f867cf3;
    ram_cell[    5209] = 32'h6cc6eb42;
    ram_cell[    5210] = 32'h35b35007;
    ram_cell[    5211] = 32'h16c77b4f;
    ram_cell[    5212] = 32'h6dc4523c;
    ram_cell[    5213] = 32'hb2f0c39d;
    ram_cell[    5214] = 32'h7558a476;
    ram_cell[    5215] = 32'hfdc92e02;
    ram_cell[    5216] = 32'h5c08140c;
    ram_cell[    5217] = 32'h02cba386;
    ram_cell[    5218] = 32'hb1d74547;
    ram_cell[    5219] = 32'heb17002f;
    ram_cell[    5220] = 32'hb1a1288e;
    ram_cell[    5221] = 32'h407838ac;
    ram_cell[    5222] = 32'h5b991c6b;
    ram_cell[    5223] = 32'h0fd378b4;
    ram_cell[    5224] = 32'hf6baa62b;
    ram_cell[    5225] = 32'hefa65e6b;
    ram_cell[    5226] = 32'hce8f4c51;
    ram_cell[    5227] = 32'h3acc4635;
    ram_cell[    5228] = 32'hf49638ad;
    ram_cell[    5229] = 32'h65c19073;
    ram_cell[    5230] = 32'h704d1c50;
    ram_cell[    5231] = 32'hbbc6e8c5;
    ram_cell[    5232] = 32'h172771e0;
    ram_cell[    5233] = 32'ha317c8a9;
    ram_cell[    5234] = 32'h1ff651e6;
    ram_cell[    5235] = 32'h3bd7a178;
    ram_cell[    5236] = 32'h1288fb30;
    ram_cell[    5237] = 32'hed746d1c;
    ram_cell[    5238] = 32'h5e1dc9e3;
    ram_cell[    5239] = 32'h80dccdf4;
    ram_cell[    5240] = 32'h70b708c9;
    ram_cell[    5241] = 32'h5101cd4f;
    ram_cell[    5242] = 32'hdffb9a6a;
    ram_cell[    5243] = 32'hafa5d5ee;
    ram_cell[    5244] = 32'hafd195ea;
    ram_cell[    5245] = 32'h71b07b5d;
    ram_cell[    5246] = 32'hf203696d;
    ram_cell[    5247] = 32'h42a4f9bd;
    ram_cell[    5248] = 32'h43ee1e00;
    ram_cell[    5249] = 32'hb0796b50;
    ram_cell[    5250] = 32'hf4609308;
    ram_cell[    5251] = 32'he6319213;
    ram_cell[    5252] = 32'h59ca8d77;
    ram_cell[    5253] = 32'hcc193672;
    ram_cell[    5254] = 32'h53e00104;
    ram_cell[    5255] = 32'h879c9349;
    ram_cell[    5256] = 32'hd468309a;
    ram_cell[    5257] = 32'he56a1a5b;
    ram_cell[    5258] = 32'h30cfe224;
    ram_cell[    5259] = 32'h37bfa4df;
    ram_cell[    5260] = 32'h825b048b;
    ram_cell[    5261] = 32'h1c082319;
    ram_cell[    5262] = 32'hf58feac7;
    ram_cell[    5263] = 32'h3db4a303;
    ram_cell[    5264] = 32'h43953380;
    ram_cell[    5265] = 32'hb12ef548;
    ram_cell[    5266] = 32'h2cb5b514;
    ram_cell[    5267] = 32'h6991823f;
    ram_cell[    5268] = 32'hc16e96ff;
    ram_cell[    5269] = 32'h7cd71e7f;
    ram_cell[    5270] = 32'hcf556152;
    ram_cell[    5271] = 32'h3e6c7988;
    ram_cell[    5272] = 32'h3d0ac382;
    ram_cell[    5273] = 32'h0b11fa8a;
    ram_cell[    5274] = 32'hb0adcc6b;
    ram_cell[    5275] = 32'h9616896f;
    ram_cell[    5276] = 32'ha5b0dcb6;
    ram_cell[    5277] = 32'h235a5f0b;
    ram_cell[    5278] = 32'hf1b13ac9;
    ram_cell[    5279] = 32'hf7e3c142;
    ram_cell[    5280] = 32'hc3941f6a;
    ram_cell[    5281] = 32'hda0fc94a;
    ram_cell[    5282] = 32'h0fc28fb7;
    ram_cell[    5283] = 32'h134694c8;
    ram_cell[    5284] = 32'h16ff22f1;
    ram_cell[    5285] = 32'h403dd2f4;
    ram_cell[    5286] = 32'ha8b34632;
    ram_cell[    5287] = 32'h62c62d3d;
    ram_cell[    5288] = 32'ha78d570c;
    ram_cell[    5289] = 32'h1c7121a8;
    ram_cell[    5290] = 32'h485b0d6d;
    ram_cell[    5291] = 32'hceec76ba;
    ram_cell[    5292] = 32'h9d6ac2ac;
    ram_cell[    5293] = 32'h6147deaa;
    ram_cell[    5294] = 32'h3b28c467;
    ram_cell[    5295] = 32'h28720108;
    ram_cell[    5296] = 32'hb84ddfd3;
    ram_cell[    5297] = 32'hae029e96;
    ram_cell[    5298] = 32'h45e85984;
    ram_cell[    5299] = 32'hc5bde766;
    ram_cell[    5300] = 32'hd675da80;
    ram_cell[    5301] = 32'he20d1b60;
    ram_cell[    5302] = 32'h7892ff0b;
    ram_cell[    5303] = 32'h780b4b90;
    ram_cell[    5304] = 32'h126eb619;
    ram_cell[    5305] = 32'h360b7c55;
    ram_cell[    5306] = 32'h8a011856;
    ram_cell[    5307] = 32'h87538a68;
    ram_cell[    5308] = 32'he55747f2;
    ram_cell[    5309] = 32'h5978284a;
    ram_cell[    5310] = 32'hc5b2105e;
    ram_cell[    5311] = 32'hcd0e5de5;
    ram_cell[    5312] = 32'h551b4221;
    ram_cell[    5313] = 32'h2ca395d8;
    ram_cell[    5314] = 32'h26979f7b;
    ram_cell[    5315] = 32'ha868680a;
    ram_cell[    5316] = 32'h876f01b2;
    ram_cell[    5317] = 32'h12de3a60;
    ram_cell[    5318] = 32'hda55eb93;
    ram_cell[    5319] = 32'h270b6310;
    ram_cell[    5320] = 32'hf8676355;
    ram_cell[    5321] = 32'h79844f63;
    ram_cell[    5322] = 32'h733ae731;
    ram_cell[    5323] = 32'h8b902391;
    ram_cell[    5324] = 32'hdeb6425b;
    ram_cell[    5325] = 32'h2dfc5104;
    ram_cell[    5326] = 32'h43435ce7;
    ram_cell[    5327] = 32'hc5e77bd5;
    ram_cell[    5328] = 32'h86346f6a;
    ram_cell[    5329] = 32'h32f3d22d;
    ram_cell[    5330] = 32'hbefb58ee;
    ram_cell[    5331] = 32'hd7fb4cd0;
    ram_cell[    5332] = 32'h0d23cdb1;
    ram_cell[    5333] = 32'hf293b020;
    ram_cell[    5334] = 32'hee2fb56d;
    ram_cell[    5335] = 32'hcedd7177;
    ram_cell[    5336] = 32'h3f770d50;
    ram_cell[    5337] = 32'hef18b633;
    ram_cell[    5338] = 32'h4a854cba;
    ram_cell[    5339] = 32'h521a0e43;
    ram_cell[    5340] = 32'h9229f399;
    ram_cell[    5341] = 32'habb03f88;
    ram_cell[    5342] = 32'h78347935;
    ram_cell[    5343] = 32'hc8773b01;
    ram_cell[    5344] = 32'he0401173;
    ram_cell[    5345] = 32'he4225945;
    ram_cell[    5346] = 32'h0a8f481a;
    ram_cell[    5347] = 32'h2c985740;
    ram_cell[    5348] = 32'h113a0157;
    ram_cell[    5349] = 32'hd7cb7197;
    ram_cell[    5350] = 32'hff70648b;
    ram_cell[    5351] = 32'hc6403acd;
    ram_cell[    5352] = 32'hb631f36a;
    ram_cell[    5353] = 32'hb4f17728;
    ram_cell[    5354] = 32'hd7761374;
    ram_cell[    5355] = 32'hf47376c6;
    ram_cell[    5356] = 32'hdfcefbeb;
    ram_cell[    5357] = 32'h783bac5e;
    ram_cell[    5358] = 32'hd291005c;
    ram_cell[    5359] = 32'hf9155e3f;
    ram_cell[    5360] = 32'hc0c0694a;
    ram_cell[    5361] = 32'hb48837d1;
    ram_cell[    5362] = 32'h0151a541;
    ram_cell[    5363] = 32'h9ec9c374;
    ram_cell[    5364] = 32'h25a79e68;
    ram_cell[    5365] = 32'h3e0fae80;
    ram_cell[    5366] = 32'h6074f8fe;
    ram_cell[    5367] = 32'hb12ded28;
    ram_cell[    5368] = 32'h10bdd875;
    ram_cell[    5369] = 32'he64bd7d6;
    ram_cell[    5370] = 32'h4f64f68c;
    ram_cell[    5371] = 32'h31e5879c;
    ram_cell[    5372] = 32'h72bf21fb;
    ram_cell[    5373] = 32'h66ea9063;
    ram_cell[    5374] = 32'h09eea060;
    ram_cell[    5375] = 32'h9ca6d332;
    ram_cell[    5376] = 32'he50148c5;
    ram_cell[    5377] = 32'h08561ddf;
    ram_cell[    5378] = 32'hc39c429f;
    ram_cell[    5379] = 32'h2ff051eb;
    ram_cell[    5380] = 32'h90d3468e;
    ram_cell[    5381] = 32'h6cbf24c7;
    ram_cell[    5382] = 32'ha22500a6;
    ram_cell[    5383] = 32'h3e6849ef;
    ram_cell[    5384] = 32'h177c081c;
    ram_cell[    5385] = 32'hcabd2f11;
    ram_cell[    5386] = 32'h182d0e87;
    ram_cell[    5387] = 32'hf5551364;
    ram_cell[    5388] = 32'h15468565;
    ram_cell[    5389] = 32'h42b67052;
    ram_cell[    5390] = 32'h1025a076;
    ram_cell[    5391] = 32'h648551af;
    ram_cell[    5392] = 32'ha3b353b7;
    ram_cell[    5393] = 32'hbfc0fda2;
    ram_cell[    5394] = 32'hd22f2e76;
    ram_cell[    5395] = 32'h12ab4645;
    ram_cell[    5396] = 32'hc3abd8b0;
    ram_cell[    5397] = 32'h45ecce21;
    ram_cell[    5398] = 32'h1f8aef54;
    ram_cell[    5399] = 32'hfa3c9dde;
    ram_cell[    5400] = 32'h20b15dae;
    ram_cell[    5401] = 32'h3bf43249;
    ram_cell[    5402] = 32'hedf408ca;
    ram_cell[    5403] = 32'hd5909379;
    ram_cell[    5404] = 32'hb0fc80bf;
    ram_cell[    5405] = 32'ha7898f81;
    ram_cell[    5406] = 32'hd201031a;
    ram_cell[    5407] = 32'h859d907e;
    ram_cell[    5408] = 32'hb81e0fa7;
    ram_cell[    5409] = 32'h08bc8b42;
    ram_cell[    5410] = 32'ha593bc6f;
    ram_cell[    5411] = 32'hbc2407d0;
    ram_cell[    5412] = 32'h0aea78c2;
    ram_cell[    5413] = 32'hdcd668b1;
    ram_cell[    5414] = 32'hee6061b2;
    ram_cell[    5415] = 32'h4b0441c4;
    ram_cell[    5416] = 32'hac8ce5ba;
    ram_cell[    5417] = 32'h2bfa7faa;
    ram_cell[    5418] = 32'hca70abbb;
    ram_cell[    5419] = 32'h23d4f19d;
    ram_cell[    5420] = 32'h8ada9dc6;
    ram_cell[    5421] = 32'ha7aa936d;
    ram_cell[    5422] = 32'hadd1feb3;
    ram_cell[    5423] = 32'hda586a2b;
    ram_cell[    5424] = 32'h3fe7231d;
    ram_cell[    5425] = 32'h56e4814c;
    ram_cell[    5426] = 32'h2c4a1e15;
    ram_cell[    5427] = 32'h9391ced1;
    ram_cell[    5428] = 32'h1e7dcb2b;
    ram_cell[    5429] = 32'ha0664bab;
    ram_cell[    5430] = 32'he831e6c6;
    ram_cell[    5431] = 32'h828de8c9;
    ram_cell[    5432] = 32'hb7a02205;
    ram_cell[    5433] = 32'h1b11ecf9;
    ram_cell[    5434] = 32'h9867a1a5;
    ram_cell[    5435] = 32'h4abbad69;
    ram_cell[    5436] = 32'h2c732364;
    ram_cell[    5437] = 32'hace13307;
    ram_cell[    5438] = 32'h3003db43;
    ram_cell[    5439] = 32'h3730f80e;
    ram_cell[    5440] = 32'hc6db0eb7;
    ram_cell[    5441] = 32'h491f9226;
    ram_cell[    5442] = 32'h38d0cd24;
    ram_cell[    5443] = 32'h4e41943c;
    ram_cell[    5444] = 32'h2ec4effd;
    ram_cell[    5445] = 32'h78fc257b;
    ram_cell[    5446] = 32'h034f791a;
    ram_cell[    5447] = 32'h688bf667;
    ram_cell[    5448] = 32'hf4a3edd4;
    ram_cell[    5449] = 32'ha241f8a6;
    ram_cell[    5450] = 32'h58d5c949;
    ram_cell[    5451] = 32'h0d3dd4fb;
    ram_cell[    5452] = 32'hd5c22e01;
    ram_cell[    5453] = 32'h99f0c9fc;
    ram_cell[    5454] = 32'hb06e6ea6;
    ram_cell[    5455] = 32'hb22a6896;
    ram_cell[    5456] = 32'h560eb497;
    ram_cell[    5457] = 32'h53867413;
    ram_cell[    5458] = 32'h01a5a4a0;
    ram_cell[    5459] = 32'h6815fd05;
    ram_cell[    5460] = 32'h354e8e38;
    ram_cell[    5461] = 32'h5b7cdefc;
    ram_cell[    5462] = 32'hb0f84de5;
    ram_cell[    5463] = 32'hb8ec7248;
    ram_cell[    5464] = 32'h4a9c8c32;
    ram_cell[    5465] = 32'h10e44cd4;
    ram_cell[    5466] = 32'h527fe8c8;
    ram_cell[    5467] = 32'hb0244c74;
    ram_cell[    5468] = 32'h5e2eb5ce;
    ram_cell[    5469] = 32'h9a0afabe;
    ram_cell[    5470] = 32'h21f1e744;
    ram_cell[    5471] = 32'h07e5b62f;
    ram_cell[    5472] = 32'hd9941dbb;
    ram_cell[    5473] = 32'h7db36d6f;
    ram_cell[    5474] = 32'h2fd880ec;
    ram_cell[    5475] = 32'h7c84eadd;
    ram_cell[    5476] = 32'h4ef468cc;
    ram_cell[    5477] = 32'h2caba46f;
    ram_cell[    5478] = 32'hf16d8ab6;
    ram_cell[    5479] = 32'h419384d5;
    ram_cell[    5480] = 32'ha5821b93;
    ram_cell[    5481] = 32'hc3fa5423;
    ram_cell[    5482] = 32'h94dca565;
    ram_cell[    5483] = 32'h0d7306f9;
    ram_cell[    5484] = 32'hdb78d653;
    ram_cell[    5485] = 32'hd01abe5d;
    ram_cell[    5486] = 32'h91d2dfe1;
    ram_cell[    5487] = 32'h16bf7a6d;
    ram_cell[    5488] = 32'h46c29f35;
    ram_cell[    5489] = 32'h158bf0ff;
    ram_cell[    5490] = 32'h330b0c59;
    ram_cell[    5491] = 32'h52e994f9;
    ram_cell[    5492] = 32'hf9e274a2;
    ram_cell[    5493] = 32'hbbc2f6cf;
    ram_cell[    5494] = 32'h3845a9d3;
    ram_cell[    5495] = 32'h0f611777;
    ram_cell[    5496] = 32'h02635b50;
    ram_cell[    5497] = 32'h23c2ecf1;
    ram_cell[    5498] = 32'h9e524862;
    ram_cell[    5499] = 32'hf8687b72;
    ram_cell[    5500] = 32'h904975ae;
    ram_cell[    5501] = 32'hb44f84e6;
    ram_cell[    5502] = 32'h8279585a;
    ram_cell[    5503] = 32'hf2bf58e5;
    ram_cell[    5504] = 32'hdf4b82ac;
    ram_cell[    5505] = 32'h1805076d;
    ram_cell[    5506] = 32'h0234e89d;
    ram_cell[    5507] = 32'h365c9ae9;
    ram_cell[    5508] = 32'he8d12390;
    ram_cell[    5509] = 32'hd2e4d983;
    ram_cell[    5510] = 32'h261da0a8;
    ram_cell[    5511] = 32'hbd07264e;
    ram_cell[    5512] = 32'h20f5f392;
    ram_cell[    5513] = 32'h007a4550;
    ram_cell[    5514] = 32'hdaac11a5;
    ram_cell[    5515] = 32'hb7fae5bd;
    ram_cell[    5516] = 32'h142c9d4e;
    ram_cell[    5517] = 32'h3a659125;
    ram_cell[    5518] = 32'h45c0e15c;
    ram_cell[    5519] = 32'hc9381676;
    ram_cell[    5520] = 32'h8abd6198;
    ram_cell[    5521] = 32'h9ba3538b;
    ram_cell[    5522] = 32'h7da563af;
    ram_cell[    5523] = 32'h8b5aa081;
    ram_cell[    5524] = 32'hb9fcfcef;
    ram_cell[    5525] = 32'hf5428bbf;
    ram_cell[    5526] = 32'hf5a21763;
    ram_cell[    5527] = 32'h15c75275;
    ram_cell[    5528] = 32'h386dc6c0;
    ram_cell[    5529] = 32'h024bc997;
    ram_cell[    5530] = 32'h19f17306;
    ram_cell[    5531] = 32'h6d7a4ffe;
    ram_cell[    5532] = 32'h31af908e;
    ram_cell[    5533] = 32'h30d0c8b3;
    ram_cell[    5534] = 32'h0d0ea03f;
    ram_cell[    5535] = 32'h0d98b096;
    ram_cell[    5536] = 32'h4f0f20b9;
    ram_cell[    5537] = 32'h8efcec62;
    ram_cell[    5538] = 32'h71c027f2;
    ram_cell[    5539] = 32'h932897a9;
    ram_cell[    5540] = 32'h58707e40;
    ram_cell[    5541] = 32'h29c404ad;
    ram_cell[    5542] = 32'hffe2f7aa;
    ram_cell[    5543] = 32'hbbf0fed1;
    ram_cell[    5544] = 32'h8fd2c085;
    ram_cell[    5545] = 32'ha68d1fcd;
    ram_cell[    5546] = 32'ha8d8ec1f;
    ram_cell[    5547] = 32'h966dac83;
    ram_cell[    5548] = 32'he003dd57;
    ram_cell[    5549] = 32'h142b667d;
    ram_cell[    5550] = 32'h59e1b74f;
    ram_cell[    5551] = 32'h3eab67c1;
    ram_cell[    5552] = 32'h349d28ea;
    ram_cell[    5553] = 32'hf1f6504e;
    ram_cell[    5554] = 32'hc8506718;
    ram_cell[    5555] = 32'h0ca73ea6;
    ram_cell[    5556] = 32'h93fd7bb4;
    ram_cell[    5557] = 32'hf5a097d4;
    ram_cell[    5558] = 32'hb1c1410c;
    ram_cell[    5559] = 32'h5f87a429;
    ram_cell[    5560] = 32'hee792c43;
    ram_cell[    5561] = 32'h7f3067a2;
    ram_cell[    5562] = 32'h7b534026;
    ram_cell[    5563] = 32'h59f61ec8;
    ram_cell[    5564] = 32'h764a907d;
    ram_cell[    5565] = 32'hf40f38cd;
    ram_cell[    5566] = 32'h24f729e5;
    ram_cell[    5567] = 32'ha392b2ce;
    ram_cell[    5568] = 32'h25a84072;
    ram_cell[    5569] = 32'h0dcbae2a;
    ram_cell[    5570] = 32'h920580e8;
    ram_cell[    5571] = 32'h5b6a6ea9;
    ram_cell[    5572] = 32'h0500a13a;
    ram_cell[    5573] = 32'h5ada8a48;
    ram_cell[    5574] = 32'hc484d37c;
    ram_cell[    5575] = 32'h18991e17;
    ram_cell[    5576] = 32'h23bed994;
    ram_cell[    5577] = 32'ha8c18b19;
    ram_cell[    5578] = 32'h16f7717c;
    ram_cell[    5579] = 32'heb90b8f4;
    ram_cell[    5580] = 32'h86857e96;
    ram_cell[    5581] = 32'h457fa5c2;
    ram_cell[    5582] = 32'hf2fec1a9;
    ram_cell[    5583] = 32'h5a62fe44;
    ram_cell[    5584] = 32'h351063db;
    ram_cell[    5585] = 32'h111dc74d;
    ram_cell[    5586] = 32'h9b5fbe61;
    ram_cell[    5587] = 32'h31c25483;
    ram_cell[    5588] = 32'h5dd8d0f3;
    ram_cell[    5589] = 32'h4ed513f4;
    ram_cell[    5590] = 32'h7163c839;
    ram_cell[    5591] = 32'hfcd9b763;
    ram_cell[    5592] = 32'hc8d0dd25;
    ram_cell[    5593] = 32'h73c28020;
    ram_cell[    5594] = 32'h678d2b59;
    ram_cell[    5595] = 32'had41af74;
    ram_cell[    5596] = 32'hf30c5ff8;
    ram_cell[    5597] = 32'he6be7e81;
    ram_cell[    5598] = 32'h8a8f2466;
    ram_cell[    5599] = 32'hd071a22b;
    ram_cell[    5600] = 32'hb404e065;
    ram_cell[    5601] = 32'hac391d7d;
    ram_cell[    5602] = 32'h2eb7686d;
    ram_cell[    5603] = 32'h1799e185;
    ram_cell[    5604] = 32'hcecaf1b4;
    ram_cell[    5605] = 32'h9f1cbb1f;
    ram_cell[    5606] = 32'he6b540dc;
    ram_cell[    5607] = 32'h06f162c4;
    ram_cell[    5608] = 32'hfd25da86;
    ram_cell[    5609] = 32'h9580a5d4;
    ram_cell[    5610] = 32'h2d0fd72e;
    ram_cell[    5611] = 32'h5e8270d2;
    ram_cell[    5612] = 32'h5a7792e9;
    ram_cell[    5613] = 32'h332c2f23;
    ram_cell[    5614] = 32'h4ecc7964;
    ram_cell[    5615] = 32'hdd87956f;
    ram_cell[    5616] = 32'hf6c314e3;
    ram_cell[    5617] = 32'h12b81c84;
    ram_cell[    5618] = 32'h2550aa9e;
    ram_cell[    5619] = 32'hd3056aeb;
    ram_cell[    5620] = 32'hbc7f8f1b;
    ram_cell[    5621] = 32'h17a342e3;
    ram_cell[    5622] = 32'h46de450c;
    ram_cell[    5623] = 32'h2f76cce2;
    ram_cell[    5624] = 32'h4c18664c;
    ram_cell[    5625] = 32'h7a31b10e;
    ram_cell[    5626] = 32'hd3b6aa35;
    ram_cell[    5627] = 32'h1453ede7;
    ram_cell[    5628] = 32'h879e6a23;
    ram_cell[    5629] = 32'h4656c66a;
    ram_cell[    5630] = 32'h49deadf9;
    ram_cell[    5631] = 32'hb4e25c19;
    ram_cell[    5632] = 32'hfdb994e3;
    ram_cell[    5633] = 32'h68886d03;
    ram_cell[    5634] = 32'ha2b09ba8;
    ram_cell[    5635] = 32'h2c8e9284;
    ram_cell[    5636] = 32'hb850b746;
    ram_cell[    5637] = 32'h3bb7fed8;
    ram_cell[    5638] = 32'h229daf6b;
    ram_cell[    5639] = 32'h0a5a810e;
    ram_cell[    5640] = 32'hcf983895;
    ram_cell[    5641] = 32'h2b655cf3;
    ram_cell[    5642] = 32'hb5ac23ab;
    ram_cell[    5643] = 32'h39efd83a;
    ram_cell[    5644] = 32'h74feff68;
    ram_cell[    5645] = 32'h759f1f70;
    ram_cell[    5646] = 32'h26b49a26;
    ram_cell[    5647] = 32'h6b3f9a96;
    ram_cell[    5648] = 32'h478a013c;
    ram_cell[    5649] = 32'h7b5f59a7;
    ram_cell[    5650] = 32'h28bbce5c;
    ram_cell[    5651] = 32'h82a9e8d6;
    ram_cell[    5652] = 32'h86fc5563;
    ram_cell[    5653] = 32'h41e4b006;
    ram_cell[    5654] = 32'he89bd46f;
    ram_cell[    5655] = 32'h0e41b345;
    ram_cell[    5656] = 32'h5fe6385b;
    ram_cell[    5657] = 32'h9db152a4;
    ram_cell[    5658] = 32'h149be4f0;
    ram_cell[    5659] = 32'h5637113c;
    ram_cell[    5660] = 32'he1d157ca;
    ram_cell[    5661] = 32'h5868f552;
    ram_cell[    5662] = 32'h0e744744;
    ram_cell[    5663] = 32'h924dc4a0;
    ram_cell[    5664] = 32'hf3cd4e59;
    ram_cell[    5665] = 32'h45456054;
    ram_cell[    5666] = 32'hd7989f1c;
    ram_cell[    5667] = 32'h85f18ab8;
    ram_cell[    5668] = 32'hadb1dd35;
    ram_cell[    5669] = 32'hd6581cbe;
    ram_cell[    5670] = 32'h5b13e04c;
    ram_cell[    5671] = 32'h81231839;
    ram_cell[    5672] = 32'h57e41fc9;
    ram_cell[    5673] = 32'hdf389369;
    ram_cell[    5674] = 32'h5b874d64;
    ram_cell[    5675] = 32'h5d173f7c;
    ram_cell[    5676] = 32'hc6686f0a;
    ram_cell[    5677] = 32'h97acba2d;
    ram_cell[    5678] = 32'h6e451749;
    ram_cell[    5679] = 32'hd3c23226;
    ram_cell[    5680] = 32'h45b4ae83;
    ram_cell[    5681] = 32'h11dd6b0a;
    ram_cell[    5682] = 32'h2db5b358;
    ram_cell[    5683] = 32'h1ce6c999;
    ram_cell[    5684] = 32'h070513e8;
    ram_cell[    5685] = 32'h2b470453;
    ram_cell[    5686] = 32'h64ffb07c;
    ram_cell[    5687] = 32'hc7c711a2;
    ram_cell[    5688] = 32'h4cec08ea;
    ram_cell[    5689] = 32'hbb53c2d0;
    ram_cell[    5690] = 32'ha6e7192a;
    ram_cell[    5691] = 32'h1555db26;
    ram_cell[    5692] = 32'hfb404897;
    ram_cell[    5693] = 32'hb8133cf9;
    ram_cell[    5694] = 32'he6238755;
    ram_cell[    5695] = 32'h89b22606;
    ram_cell[    5696] = 32'hdf5fbfbe;
    ram_cell[    5697] = 32'hc4c91958;
    ram_cell[    5698] = 32'h366f2cc0;
    ram_cell[    5699] = 32'h35ec3dbe;
    ram_cell[    5700] = 32'he6031c2b;
    ram_cell[    5701] = 32'h9f762d96;
    ram_cell[    5702] = 32'h57f9c9df;
    ram_cell[    5703] = 32'h884fb591;
    ram_cell[    5704] = 32'hcc033278;
    ram_cell[    5705] = 32'h4fb592f8;
    ram_cell[    5706] = 32'ha6be3797;
    ram_cell[    5707] = 32'h6ec0d5a8;
    ram_cell[    5708] = 32'h12ed05a1;
    ram_cell[    5709] = 32'hedba6a07;
    ram_cell[    5710] = 32'h9ad42262;
    ram_cell[    5711] = 32'h3d5e0b3c;
    ram_cell[    5712] = 32'h7583470e;
    ram_cell[    5713] = 32'ha50dba51;
    ram_cell[    5714] = 32'h435852ee;
    ram_cell[    5715] = 32'h0cfd2ac5;
    ram_cell[    5716] = 32'he9fc302d;
    ram_cell[    5717] = 32'h691ad6ff;
    ram_cell[    5718] = 32'h36801299;
    ram_cell[    5719] = 32'hcf639526;
    ram_cell[    5720] = 32'h9329f4aa;
    ram_cell[    5721] = 32'hbbb73545;
    ram_cell[    5722] = 32'h4e482f82;
    ram_cell[    5723] = 32'h4d5ec17b;
    ram_cell[    5724] = 32'hb13a2e6c;
    ram_cell[    5725] = 32'hb8f00eb2;
    ram_cell[    5726] = 32'h1170ff83;
    ram_cell[    5727] = 32'hc81d1db4;
    ram_cell[    5728] = 32'hb3dd8cf7;
    ram_cell[    5729] = 32'h7072b2ca;
    ram_cell[    5730] = 32'h4e703083;
    ram_cell[    5731] = 32'hbe78bd64;
    ram_cell[    5732] = 32'h0f4b47fc;
    ram_cell[    5733] = 32'hd85a7520;
    ram_cell[    5734] = 32'hfc504d39;
    ram_cell[    5735] = 32'hfee5cbb6;
    ram_cell[    5736] = 32'hfb594f64;
    ram_cell[    5737] = 32'h18f8d889;
    ram_cell[    5738] = 32'hcc3c460d;
    ram_cell[    5739] = 32'h8852db6d;
    ram_cell[    5740] = 32'hb95597be;
    ram_cell[    5741] = 32'h35baef83;
    ram_cell[    5742] = 32'hbbf02672;
    ram_cell[    5743] = 32'h43ee8acf;
    ram_cell[    5744] = 32'hdc7a3c0e;
    ram_cell[    5745] = 32'h20096c71;
    ram_cell[    5746] = 32'hf97d70ea;
    ram_cell[    5747] = 32'hd148ad78;
    ram_cell[    5748] = 32'hdd535cd7;
    ram_cell[    5749] = 32'h11cb8bbf;
    ram_cell[    5750] = 32'h47159eef;
    ram_cell[    5751] = 32'h025beca5;
    ram_cell[    5752] = 32'h810abdd1;
    ram_cell[    5753] = 32'he476d91a;
    ram_cell[    5754] = 32'h965fbf6d;
    ram_cell[    5755] = 32'h2a4750b2;
    ram_cell[    5756] = 32'hbe0c64a8;
    ram_cell[    5757] = 32'h24a9195c;
    ram_cell[    5758] = 32'hde0ab1b2;
    ram_cell[    5759] = 32'h5acb9ba9;
    ram_cell[    5760] = 32'h95576dd7;
    ram_cell[    5761] = 32'h53e8f5ab;
    ram_cell[    5762] = 32'hdd23e0cc;
    ram_cell[    5763] = 32'h7eff5899;
    ram_cell[    5764] = 32'h65cec82d;
    ram_cell[    5765] = 32'h07eb529a;
    ram_cell[    5766] = 32'ha333d963;
    ram_cell[    5767] = 32'h42f73a8e;
    ram_cell[    5768] = 32'hae0e8d20;
    ram_cell[    5769] = 32'hec61c385;
    ram_cell[    5770] = 32'h5e39e5a8;
    ram_cell[    5771] = 32'h3f59eae3;
    ram_cell[    5772] = 32'hc09ae1ec;
    ram_cell[    5773] = 32'h9aed14bc;
    ram_cell[    5774] = 32'h8524b4fd;
    ram_cell[    5775] = 32'h564795f3;
    ram_cell[    5776] = 32'hc144f95d;
    ram_cell[    5777] = 32'h77a28bc8;
    ram_cell[    5778] = 32'h30b05941;
    ram_cell[    5779] = 32'h4d5cf2ac;
    ram_cell[    5780] = 32'h22d86bc5;
    ram_cell[    5781] = 32'hfd8bf133;
    ram_cell[    5782] = 32'h9b1ff0df;
    ram_cell[    5783] = 32'hc1476b1d;
    ram_cell[    5784] = 32'h882692a9;
    ram_cell[    5785] = 32'h481ce350;
    ram_cell[    5786] = 32'hf1841e51;
    ram_cell[    5787] = 32'hb3e49e86;
    ram_cell[    5788] = 32'h45a5be56;
    ram_cell[    5789] = 32'h80d1c5cf;
    ram_cell[    5790] = 32'hbc285258;
    ram_cell[    5791] = 32'h7addef8a;
    ram_cell[    5792] = 32'h497411bc;
    ram_cell[    5793] = 32'h20975eb7;
    ram_cell[    5794] = 32'h57662e9e;
    ram_cell[    5795] = 32'ha9a6b6fe;
    ram_cell[    5796] = 32'h56dc8acf;
    ram_cell[    5797] = 32'h2252019d;
    ram_cell[    5798] = 32'h5119d288;
    ram_cell[    5799] = 32'h1fd2dc68;
    ram_cell[    5800] = 32'h57cbbe28;
    ram_cell[    5801] = 32'h4286270e;
    ram_cell[    5802] = 32'hf05f2ce3;
    ram_cell[    5803] = 32'h7249fc37;
    ram_cell[    5804] = 32'hb4b3c3dc;
    ram_cell[    5805] = 32'hd46ee39d;
    ram_cell[    5806] = 32'h14e68465;
    ram_cell[    5807] = 32'h1233041b;
    ram_cell[    5808] = 32'h2c2a20f0;
    ram_cell[    5809] = 32'hb3a0a37b;
    ram_cell[    5810] = 32'h3ccb62a3;
    ram_cell[    5811] = 32'h2abf8f5c;
    ram_cell[    5812] = 32'h4b9339d4;
    ram_cell[    5813] = 32'h64aa606d;
    ram_cell[    5814] = 32'hcc119f9f;
    ram_cell[    5815] = 32'hf0aef426;
    ram_cell[    5816] = 32'h67cdb5ac;
    ram_cell[    5817] = 32'hb2547501;
    ram_cell[    5818] = 32'hb73cb641;
    ram_cell[    5819] = 32'h1cd32e0e;
    ram_cell[    5820] = 32'he0b5d029;
    ram_cell[    5821] = 32'h322eaecf;
    ram_cell[    5822] = 32'h4385456e;
    ram_cell[    5823] = 32'h6d78fbb3;
    ram_cell[    5824] = 32'hcb45fb4a;
    ram_cell[    5825] = 32'h2483f369;
    ram_cell[    5826] = 32'he76f9b61;
    ram_cell[    5827] = 32'hb759bd3b;
    ram_cell[    5828] = 32'h88b77828;
    ram_cell[    5829] = 32'h66db82ee;
    ram_cell[    5830] = 32'h3437c331;
    ram_cell[    5831] = 32'h17b22a88;
    ram_cell[    5832] = 32'h2f72c98d;
    ram_cell[    5833] = 32'he71f87ea;
    ram_cell[    5834] = 32'hd9a9de99;
    ram_cell[    5835] = 32'hf17bba35;
    ram_cell[    5836] = 32'h32525300;
    ram_cell[    5837] = 32'hf65e047a;
    ram_cell[    5838] = 32'h59ab9ec3;
    ram_cell[    5839] = 32'h9c28d77f;
    ram_cell[    5840] = 32'h584a1682;
    ram_cell[    5841] = 32'he4d5883e;
    ram_cell[    5842] = 32'h8cc57986;
    ram_cell[    5843] = 32'h189d83db;
    ram_cell[    5844] = 32'h41f5e714;
    ram_cell[    5845] = 32'hdd3a7a0c;
    ram_cell[    5846] = 32'h6ab2c870;
    ram_cell[    5847] = 32'h7a0ef825;
    ram_cell[    5848] = 32'hc2302ab4;
    ram_cell[    5849] = 32'h9545fd7e;
    ram_cell[    5850] = 32'h4ab33387;
    ram_cell[    5851] = 32'h67324e1b;
    ram_cell[    5852] = 32'h2f2d815d;
    ram_cell[    5853] = 32'h332c8e01;
    ram_cell[    5854] = 32'he6954f9b;
    ram_cell[    5855] = 32'h73cfc854;
    ram_cell[    5856] = 32'h5fcf75a7;
    ram_cell[    5857] = 32'h1a9a6fab;
    ram_cell[    5858] = 32'h3b87c9dd;
    ram_cell[    5859] = 32'h17ce9bec;
    ram_cell[    5860] = 32'h4ad9b5db;
    ram_cell[    5861] = 32'hb7bf3cfd;
    ram_cell[    5862] = 32'he223f2bb;
    ram_cell[    5863] = 32'hc89f07fe;
    ram_cell[    5864] = 32'h4794f386;
    ram_cell[    5865] = 32'h7c049184;
    ram_cell[    5866] = 32'h8f486687;
    ram_cell[    5867] = 32'hfc041284;
    ram_cell[    5868] = 32'hb9ab8c87;
    ram_cell[    5869] = 32'hd1c8a7f5;
    ram_cell[    5870] = 32'h5b254b0e;
    ram_cell[    5871] = 32'hc3b59885;
    ram_cell[    5872] = 32'hb1b54f64;
    ram_cell[    5873] = 32'he2cf0ce9;
    ram_cell[    5874] = 32'h71dd4a66;
    ram_cell[    5875] = 32'ha46d5052;
    ram_cell[    5876] = 32'h9a67ff91;
    ram_cell[    5877] = 32'h8175072c;
    ram_cell[    5878] = 32'h037bb24d;
    ram_cell[    5879] = 32'hf5b61507;
    ram_cell[    5880] = 32'hf86dc7ac;
    ram_cell[    5881] = 32'h5c8e63d0;
    ram_cell[    5882] = 32'h035a5fd1;
    ram_cell[    5883] = 32'h8a5f7535;
    ram_cell[    5884] = 32'h87001062;
    ram_cell[    5885] = 32'h63d7763f;
    ram_cell[    5886] = 32'h26ea9214;
    ram_cell[    5887] = 32'h86c06ef1;
    ram_cell[    5888] = 32'h77025f14;
    ram_cell[    5889] = 32'hd7626ed6;
    ram_cell[    5890] = 32'h5faf1f15;
    ram_cell[    5891] = 32'hfcdc0138;
    ram_cell[    5892] = 32'hcc3df038;
    ram_cell[    5893] = 32'hf081ac24;
    ram_cell[    5894] = 32'hb5a9d0a6;
    ram_cell[    5895] = 32'h02c76c1a;
    ram_cell[    5896] = 32'h0454cd83;
    ram_cell[    5897] = 32'h40c831f0;
    ram_cell[    5898] = 32'hba609d96;
    ram_cell[    5899] = 32'he6a61e3e;
    ram_cell[    5900] = 32'h6eb5c770;
    ram_cell[    5901] = 32'h05d42abe;
    ram_cell[    5902] = 32'hc1baf1f9;
    ram_cell[    5903] = 32'h27239627;
    ram_cell[    5904] = 32'he10b6b2d;
    ram_cell[    5905] = 32'h712fabb8;
    ram_cell[    5906] = 32'h28060aa5;
    ram_cell[    5907] = 32'hb32d9621;
    ram_cell[    5908] = 32'h212b086e;
    ram_cell[    5909] = 32'h5e603870;
    ram_cell[    5910] = 32'h46ab414a;
    ram_cell[    5911] = 32'h7fa1434e;
    ram_cell[    5912] = 32'h59eee21a;
    ram_cell[    5913] = 32'h67a27ea6;
    ram_cell[    5914] = 32'h55b5fc49;
    ram_cell[    5915] = 32'h43710f7c;
    ram_cell[    5916] = 32'hc37cd5f5;
    ram_cell[    5917] = 32'h1d305136;
    ram_cell[    5918] = 32'h3fe9eafb;
    ram_cell[    5919] = 32'hfffe8576;
    ram_cell[    5920] = 32'hb2b3e511;
    ram_cell[    5921] = 32'ha0b36e45;
    ram_cell[    5922] = 32'hc537c97c;
    ram_cell[    5923] = 32'h4a5d8290;
    ram_cell[    5924] = 32'hf95c6602;
    ram_cell[    5925] = 32'h365e23cf;
    ram_cell[    5926] = 32'hc5012289;
    ram_cell[    5927] = 32'h840b5f87;
    ram_cell[    5928] = 32'hc4ea790b;
    ram_cell[    5929] = 32'he46cf4dc;
    ram_cell[    5930] = 32'ha3134c3e;
    ram_cell[    5931] = 32'hc7f71248;
    ram_cell[    5932] = 32'h27cd24d6;
    ram_cell[    5933] = 32'h221967c9;
    ram_cell[    5934] = 32'hd5653b1a;
    ram_cell[    5935] = 32'h49e662f8;
    ram_cell[    5936] = 32'hdd4add3f;
    ram_cell[    5937] = 32'h0d3f2f85;
    ram_cell[    5938] = 32'hb87dbb03;
    ram_cell[    5939] = 32'h15aa6770;
    ram_cell[    5940] = 32'hd25fac05;
    ram_cell[    5941] = 32'h3d509f93;
    ram_cell[    5942] = 32'h870f8585;
    ram_cell[    5943] = 32'hdc488411;
    ram_cell[    5944] = 32'h16b621d0;
    ram_cell[    5945] = 32'hfd5acb48;
    ram_cell[    5946] = 32'ha6475dd2;
    ram_cell[    5947] = 32'h26c41980;
    ram_cell[    5948] = 32'h33bd63d1;
    ram_cell[    5949] = 32'h5555b3c0;
    ram_cell[    5950] = 32'h0548b32c;
    ram_cell[    5951] = 32'hb35f17dc;
    ram_cell[    5952] = 32'h3b60f9b5;
    ram_cell[    5953] = 32'h45ccf335;
    ram_cell[    5954] = 32'h8b906971;
    ram_cell[    5955] = 32'h37a94b22;
    ram_cell[    5956] = 32'h051c6ab5;
    ram_cell[    5957] = 32'he83a3f51;
    ram_cell[    5958] = 32'h934a6b14;
    ram_cell[    5959] = 32'hbbd62581;
    ram_cell[    5960] = 32'hc402cfc4;
    ram_cell[    5961] = 32'hd4a7bdbb;
    ram_cell[    5962] = 32'hdd9837fa;
    ram_cell[    5963] = 32'h3c3573bf;
    ram_cell[    5964] = 32'h34ece145;
    ram_cell[    5965] = 32'hdde6622b;
    ram_cell[    5966] = 32'hebb4e925;
    ram_cell[    5967] = 32'h89bdac6d;
    ram_cell[    5968] = 32'hac49a19e;
    ram_cell[    5969] = 32'h071ab90a;
    ram_cell[    5970] = 32'hc70c2148;
    ram_cell[    5971] = 32'h569c502d;
    ram_cell[    5972] = 32'h2c32f9ab;
    ram_cell[    5973] = 32'h9ba6f91e;
    ram_cell[    5974] = 32'h9b4345f7;
    ram_cell[    5975] = 32'hff729ecf;
    ram_cell[    5976] = 32'h939ffe8a;
    ram_cell[    5977] = 32'h71d1f3cf;
    ram_cell[    5978] = 32'h32f1e886;
    ram_cell[    5979] = 32'hbe6dbcab;
    ram_cell[    5980] = 32'h18f534e1;
    ram_cell[    5981] = 32'he7df48b5;
    ram_cell[    5982] = 32'h60adb046;
    ram_cell[    5983] = 32'h8bb66584;
    ram_cell[    5984] = 32'h416607b9;
    ram_cell[    5985] = 32'hb399ea06;
    ram_cell[    5986] = 32'h8c668115;
    ram_cell[    5987] = 32'h2589a7e3;
    ram_cell[    5988] = 32'h54188b56;
    ram_cell[    5989] = 32'h6870f394;
    ram_cell[    5990] = 32'ha7672cda;
    ram_cell[    5991] = 32'h52f5e948;
    ram_cell[    5992] = 32'hb511930e;
    ram_cell[    5993] = 32'hba7addd7;
    ram_cell[    5994] = 32'hd1c97c12;
    ram_cell[    5995] = 32'he42bdb45;
    ram_cell[    5996] = 32'h97157734;
    ram_cell[    5997] = 32'hbca9a29d;
    ram_cell[    5998] = 32'hfdcbeeaf;
    ram_cell[    5999] = 32'h5cefd35b;
    ram_cell[    6000] = 32'h95684512;
    ram_cell[    6001] = 32'hd446fbac;
    ram_cell[    6002] = 32'h7425c39f;
    ram_cell[    6003] = 32'h444c7ce6;
    ram_cell[    6004] = 32'hf8c8ac8a;
    ram_cell[    6005] = 32'hf6d180fe;
    ram_cell[    6006] = 32'h08c5313f;
    ram_cell[    6007] = 32'h3cbfc025;
    ram_cell[    6008] = 32'hf647b32c;
    ram_cell[    6009] = 32'ha59227d5;
    ram_cell[    6010] = 32'h556c1c82;
    ram_cell[    6011] = 32'h17039789;
    ram_cell[    6012] = 32'h1df6cbfe;
    ram_cell[    6013] = 32'h4ab65fa2;
    ram_cell[    6014] = 32'h29672800;
    ram_cell[    6015] = 32'h8106380f;
    ram_cell[    6016] = 32'hc3505f51;
    ram_cell[    6017] = 32'h812ddd39;
    ram_cell[    6018] = 32'hb0f9195c;
    ram_cell[    6019] = 32'h9d66e35d;
    ram_cell[    6020] = 32'hb0adffda;
    ram_cell[    6021] = 32'hccd3cf44;
    ram_cell[    6022] = 32'h23a3558c;
    ram_cell[    6023] = 32'h8ca4c936;
    ram_cell[    6024] = 32'h70ea5828;
    ram_cell[    6025] = 32'h7d4bcdc1;
    ram_cell[    6026] = 32'hecdc471a;
    ram_cell[    6027] = 32'hdd56b904;
    ram_cell[    6028] = 32'hc902bd47;
    ram_cell[    6029] = 32'h2193494a;
    ram_cell[    6030] = 32'ha30b439d;
    ram_cell[    6031] = 32'h57460c1a;
    ram_cell[    6032] = 32'h05c0887f;
    ram_cell[    6033] = 32'h7bfa292b;
    ram_cell[    6034] = 32'h9164e737;
    ram_cell[    6035] = 32'h4a396833;
    ram_cell[    6036] = 32'h8de0f9a9;
    ram_cell[    6037] = 32'h3cbb66a6;
    ram_cell[    6038] = 32'hfff2bf4f;
    ram_cell[    6039] = 32'hf2dce007;
    ram_cell[    6040] = 32'ha8e96f65;
    ram_cell[    6041] = 32'ha7ec5084;
    ram_cell[    6042] = 32'h327d7c13;
    ram_cell[    6043] = 32'h1380fc38;
    ram_cell[    6044] = 32'h25c8c398;
    ram_cell[    6045] = 32'h1a0843fd;
    ram_cell[    6046] = 32'hf98a8a60;
    ram_cell[    6047] = 32'hbbf3ff6c;
    ram_cell[    6048] = 32'hc50dad55;
    ram_cell[    6049] = 32'hd8833b07;
    ram_cell[    6050] = 32'h76864c5b;
    ram_cell[    6051] = 32'h907cd15e;
    ram_cell[    6052] = 32'h4be72d4a;
    ram_cell[    6053] = 32'h723bcc5e;
    ram_cell[    6054] = 32'hb10d1034;
    ram_cell[    6055] = 32'h4f1422ef;
    ram_cell[    6056] = 32'ha88b6d03;
    ram_cell[    6057] = 32'h5ad103bc;
    ram_cell[    6058] = 32'h9dc8548b;
    ram_cell[    6059] = 32'hf28d85fe;
    ram_cell[    6060] = 32'h91983dcf;
    ram_cell[    6061] = 32'h6b6dab35;
    ram_cell[    6062] = 32'hfbe2b705;
    ram_cell[    6063] = 32'hcbd2ca58;
    ram_cell[    6064] = 32'hc4458577;
    ram_cell[    6065] = 32'hcd56cc95;
    ram_cell[    6066] = 32'h1d0e0492;
    ram_cell[    6067] = 32'hef48ccf2;
    ram_cell[    6068] = 32'hb1d1f403;
    ram_cell[    6069] = 32'hb6330fa4;
    ram_cell[    6070] = 32'hd4deb7d5;
    ram_cell[    6071] = 32'h094f1afa;
    ram_cell[    6072] = 32'ha60a0c5b;
    ram_cell[    6073] = 32'hc03acb67;
    ram_cell[    6074] = 32'he7dd9308;
    ram_cell[    6075] = 32'hc73eef6b;
    ram_cell[    6076] = 32'hef434578;
    ram_cell[    6077] = 32'h40078d37;
    ram_cell[    6078] = 32'h414c48ef;
    ram_cell[    6079] = 32'h677ad857;
    ram_cell[    6080] = 32'hda9a5ee1;
    ram_cell[    6081] = 32'hcf854c86;
    ram_cell[    6082] = 32'h408a8861;
    ram_cell[    6083] = 32'h442c8f32;
    ram_cell[    6084] = 32'h2485775b;
    ram_cell[    6085] = 32'h2cd2ff1a;
    ram_cell[    6086] = 32'h6735ceff;
    ram_cell[    6087] = 32'h62b43f78;
    ram_cell[    6088] = 32'h5fd07dcd;
    ram_cell[    6089] = 32'h6666dc2d;
    ram_cell[    6090] = 32'h7094e075;
    ram_cell[    6091] = 32'hcac25d5b;
    ram_cell[    6092] = 32'h95231153;
    ram_cell[    6093] = 32'hcd244481;
    ram_cell[    6094] = 32'h345ad515;
    ram_cell[    6095] = 32'h00389585;
    ram_cell[    6096] = 32'h19310ee1;
    ram_cell[    6097] = 32'h24f7a49c;
    ram_cell[    6098] = 32'h50b4d5ca;
    ram_cell[    6099] = 32'h20d04d61;
    ram_cell[    6100] = 32'hd98fdfd1;
    ram_cell[    6101] = 32'h2692292b;
    ram_cell[    6102] = 32'h6affd5da;
    ram_cell[    6103] = 32'hd63f6017;
    ram_cell[    6104] = 32'hd922aa99;
    ram_cell[    6105] = 32'h4a9a7d96;
    ram_cell[    6106] = 32'h98215bca;
    ram_cell[    6107] = 32'h3453dc1a;
    ram_cell[    6108] = 32'hb5a5cca1;
    ram_cell[    6109] = 32'hc5e5b3d2;
    ram_cell[    6110] = 32'h6fc69bf7;
    ram_cell[    6111] = 32'hd5ead7c2;
    ram_cell[    6112] = 32'h1ca6aece;
    ram_cell[    6113] = 32'h16fe2be1;
    ram_cell[    6114] = 32'h3d12ea45;
    ram_cell[    6115] = 32'hbbf45538;
    ram_cell[    6116] = 32'h53a753f8;
    ram_cell[    6117] = 32'h5807dda6;
    ram_cell[    6118] = 32'hce044b23;
    ram_cell[    6119] = 32'h8d340206;
    ram_cell[    6120] = 32'h27aa1ad7;
    ram_cell[    6121] = 32'h8e55b967;
    ram_cell[    6122] = 32'hd3d6b6e1;
    ram_cell[    6123] = 32'h69162da1;
    ram_cell[    6124] = 32'he8177b6a;
    ram_cell[    6125] = 32'h309b9d93;
    ram_cell[    6126] = 32'hfa176ba2;
    ram_cell[    6127] = 32'h9408cddd;
    ram_cell[    6128] = 32'hd726cb2b;
    ram_cell[    6129] = 32'hb96e6fad;
    ram_cell[    6130] = 32'h4d7af38a;
    ram_cell[    6131] = 32'hb75fd097;
    ram_cell[    6132] = 32'ha5e499af;
    ram_cell[    6133] = 32'h134e28d6;
    ram_cell[    6134] = 32'hf7d904e9;
    ram_cell[    6135] = 32'hc7fd6406;
    ram_cell[    6136] = 32'h299b2a7a;
    ram_cell[    6137] = 32'hc06b38fe;
    ram_cell[    6138] = 32'h78998966;
    ram_cell[    6139] = 32'h9f7011fa;
    ram_cell[    6140] = 32'h569f6f60;
    ram_cell[    6141] = 32'h79e312eb;
    ram_cell[    6142] = 32'h7ebe15c1;
    ram_cell[    6143] = 32'hfb18bc2b;
    ram_cell[    6144] = 32'hf3b0214a;
    ram_cell[    6145] = 32'h89d80581;
    ram_cell[    6146] = 32'he0fdedba;
    ram_cell[    6147] = 32'hf285bd07;
    ram_cell[    6148] = 32'hc684d6c1;
    ram_cell[    6149] = 32'h25cfdc1e;
    ram_cell[    6150] = 32'h01e02623;
    ram_cell[    6151] = 32'hc1cc01c4;
    ram_cell[    6152] = 32'h7bda6704;
    ram_cell[    6153] = 32'h7cbee725;
    ram_cell[    6154] = 32'h533bf9aa;
    ram_cell[    6155] = 32'h3aee7186;
    ram_cell[    6156] = 32'h0f0397d0;
    ram_cell[    6157] = 32'hf0481cdb;
    ram_cell[    6158] = 32'hd18f0f34;
    ram_cell[    6159] = 32'h6fb24bcd;
    ram_cell[    6160] = 32'h41a8fd12;
    ram_cell[    6161] = 32'h188fef2c;
    ram_cell[    6162] = 32'hc04074c6;
    ram_cell[    6163] = 32'h4db6d9e2;
    ram_cell[    6164] = 32'h56ecc381;
    ram_cell[    6165] = 32'hc719909f;
    ram_cell[    6166] = 32'h3d557c21;
    ram_cell[    6167] = 32'hddfb060f;
    ram_cell[    6168] = 32'h95cf5cf0;
    ram_cell[    6169] = 32'h3c19f953;
    ram_cell[    6170] = 32'h3a10eaba;
    ram_cell[    6171] = 32'hb16e454a;
    ram_cell[    6172] = 32'h26b93d71;
    ram_cell[    6173] = 32'h4e354e01;
    ram_cell[    6174] = 32'h160e637c;
    ram_cell[    6175] = 32'h5d49af14;
    ram_cell[    6176] = 32'h814ab88b;
    ram_cell[    6177] = 32'ha3c93bcd;
    ram_cell[    6178] = 32'h9173ab16;
    ram_cell[    6179] = 32'h4bc38c07;
    ram_cell[    6180] = 32'hf25f8b7b;
    ram_cell[    6181] = 32'h25186824;
    ram_cell[    6182] = 32'h9e03cff3;
    ram_cell[    6183] = 32'he4459b45;
    ram_cell[    6184] = 32'he606a49d;
    ram_cell[    6185] = 32'h2eda1776;
    ram_cell[    6186] = 32'hb4d3a7ed;
    ram_cell[    6187] = 32'hd3ff22fe;
    ram_cell[    6188] = 32'hade10fdf;
    ram_cell[    6189] = 32'hb0f50bc6;
    ram_cell[    6190] = 32'hcc9bd23a;
    ram_cell[    6191] = 32'h81760006;
    ram_cell[    6192] = 32'h835547d5;
    ram_cell[    6193] = 32'h114cd5ae;
    ram_cell[    6194] = 32'h2b80153b;
    ram_cell[    6195] = 32'hc6851d84;
    ram_cell[    6196] = 32'h4d5d7ac4;
    ram_cell[    6197] = 32'hf144e041;
    ram_cell[    6198] = 32'h7e434d75;
    ram_cell[    6199] = 32'h8fc8f182;
    ram_cell[    6200] = 32'h209f749d;
    ram_cell[    6201] = 32'h3afeabb4;
    ram_cell[    6202] = 32'h67c0aacd;
    ram_cell[    6203] = 32'ha1511849;
    ram_cell[    6204] = 32'hce543f7f;
    ram_cell[    6205] = 32'h5bac1c13;
    ram_cell[    6206] = 32'h39cc49f9;
    ram_cell[    6207] = 32'hf2463579;
    ram_cell[    6208] = 32'he91eb2ac;
    ram_cell[    6209] = 32'hb0e93f85;
    ram_cell[    6210] = 32'h7a32f137;
    ram_cell[    6211] = 32'h4b938000;
    ram_cell[    6212] = 32'hcc0e32eb;
    ram_cell[    6213] = 32'hf9d51071;
    ram_cell[    6214] = 32'h8247c9b8;
    ram_cell[    6215] = 32'h9a8567ec;
    ram_cell[    6216] = 32'h324f0d15;
    ram_cell[    6217] = 32'h231bda45;
    ram_cell[    6218] = 32'hde1454a7;
    ram_cell[    6219] = 32'h77472ed1;
    ram_cell[    6220] = 32'h8308b091;
    ram_cell[    6221] = 32'h46172865;
    ram_cell[    6222] = 32'hfea1acb3;
    ram_cell[    6223] = 32'h0c13990c;
    ram_cell[    6224] = 32'h652a1305;
    ram_cell[    6225] = 32'h4f9b57b5;
    ram_cell[    6226] = 32'hbcf3d341;
    ram_cell[    6227] = 32'h9e6a4656;
    ram_cell[    6228] = 32'h232639f3;
    ram_cell[    6229] = 32'h01674725;
    ram_cell[    6230] = 32'hc830ffc8;
    ram_cell[    6231] = 32'h162edcbe;
    ram_cell[    6232] = 32'h44a51bad;
    ram_cell[    6233] = 32'h9080f100;
    ram_cell[    6234] = 32'he0b0fe24;
    ram_cell[    6235] = 32'h6a8c2f26;
    ram_cell[    6236] = 32'he7f65b4f;
    ram_cell[    6237] = 32'h90b19937;
    ram_cell[    6238] = 32'hdbdb80cc;
    ram_cell[    6239] = 32'h2e3c2e11;
    ram_cell[    6240] = 32'hac42c59e;
    ram_cell[    6241] = 32'h19419ce3;
    ram_cell[    6242] = 32'he1536564;
    ram_cell[    6243] = 32'hd0708e14;
    ram_cell[    6244] = 32'h305a5325;
    ram_cell[    6245] = 32'hbf82f3f1;
    ram_cell[    6246] = 32'h95718fd5;
    ram_cell[    6247] = 32'hfca73676;
    ram_cell[    6248] = 32'h90275283;
    ram_cell[    6249] = 32'hd1af9300;
    ram_cell[    6250] = 32'h8b682cbe;
    ram_cell[    6251] = 32'he8c25dea;
    ram_cell[    6252] = 32'h2101b2d3;
    ram_cell[    6253] = 32'h20c6ad39;
    ram_cell[    6254] = 32'hb5b2aa01;
    ram_cell[    6255] = 32'h8c91018c;
    ram_cell[    6256] = 32'ha33bb1a3;
    ram_cell[    6257] = 32'hbf3df0eb;
    ram_cell[    6258] = 32'ha6492e3e;
    ram_cell[    6259] = 32'hc7a85d6c;
    ram_cell[    6260] = 32'he5954c50;
    ram_cell[    6261] = 32'he50038ea;
    ram_cell[    6262] = 32'hdbca28ea;
    ram_cell[    6263] = 32'h65f98b79;
    ram_cell[    6264] = 32'h69ee9a41;
    ram_cell[    6265] = 32'ha90fbe59;
    ram_cell[    6266] = 32'h6f031365;
    ram_cell[    6267] = 32'h127ab65d;
    ram_cell[    6268] = 32'h012d84ac;
    ram_cell[    6269] = 32'h62605c1e;
    ram_cell[    6270] = 32'h90923893;
    ram_cell[    6271] = 32'hc2a9790a;
    ram_cell[    6272] = 32'h47ed23f9;
    ram_cell[    6273] = 32'hb30e99f4;
    ram_cell[    6274] = 32'hb69f6285;
    ram_cell[    6275] = 32'hb4bc0c07;
    ram_cell[    6276] = 32'h2042fedf;
    ram_cell[    6277] = 32'hb51507ce;
    ram_cell[    6278] = 32'h3e92a5a8;
    ram_cell[    6279] = 32'h3ef56488;
    ram_cell[    6280] = 32'hd0ef0e8f;
    ram_cell[    6281] = 32'h6193d1da;
    ram_cell[    6282] = 32'h361b94b0;
    ram_cell[    6283] = 32'h403fa70c;
    ram_cell[    6284] = 32'hf489ef98;
    ram_cell[    6285] = 32'h502bdbb8;
    ram_cell[    6286] = 32'h45d4b40f;
    ram_cell[    6287] = 32'h3db417a9;
    ram_cell[    6288] = 32'h6992c828;
    ram_cell[    6289] = 32'h9bf72a0b;
    ram_cell[    6290] = 32'h3d474507;
    ram_cell[    6291] = 32'ha9efec43;
    ram_cell[    6292] = 32'hf7109912;
    ram_cell[    6293] = 32'hdc296786;
    ram_cell[    6294] = 32'hc6981d7f;
    ram_cell[    6295] = 32'hc8074a77;
    ram_cell[    6296] = 32'h90d0ddae;
    ram_cell[    6297] = 32'h25f3d54a;
    ram_cell[    6298] = 32'h337980ea;
    ram_cell[    6299] = 32'h45d2bd09;
    ram_cell[    6300] = 32'hbd3a0984;
    ram_cell[    6301] = 32'h8e67a715;
    ram_cell[    6302] = 32'hffe557fc;
    ram_cell[    6303] = 32'haa556047;
    ram_cell[    6304] = 32'hea85b490;
    ram_cell[    6305] = 32'h82cc4562;
    ram_cell[    6306] = 32'hf0fb7260;
    ram_cell[    6307] = 32'h37208e75;
    ram_cell[    6308] = 32'h3ac1f100;
    ram_cell[    6309] = 32'hab70e2b8;
    ram_cell[    6310] = 32'hdf43111c;
    ram_cell[    6311] = 32'hafdf20e4;
    ram_cell[    6312] = 32'hc40af49b;
    ram_cell[    6313] = 32'h09d04a4b;
    ram_cell[    6314] = 32'h114273e5;
    ram_cell[    6315] = 32'h9295acde;
    ram_cell[    6316] = 32'h1030f48b;
    ram_cell[    6317] = 32'h3b475e9a;
    ram_cell[    6318] = 32'hddee6850;
    ram_cell[    6319] = 32'h891d22b4;
    ram_cell[    6320] = 32'hc2bee74d;
    ram_cell[    6321] = 32'h0483b6f7;
    ram_cell[    6322] = 32'h0fa07e04;
    ram_cell[    6323] = 32'h353bc263;
    ram_cell[    6324] = 32'hf2c0d386;
    ram_cell[    6325] = 32'h53cd8933;
    ram_cell[    6326] = 32'hf42b835d;
    ram_cell[    6327] = 32'h179e2a1f;
    ram_cell[    6328] = 32'h6a1ab1f2;
    ram_cell[    6329] = 32'h8d92949f;
    ram_cell[    6330] = 32'h7f858745;
    ram_cell[    6331] = 32'h1ca6d54f;
    ram_cell[    6332] = 32'h2e7ecd8a;
    ram_cell[    6333] = 32'h9e1523d3;
    ram_cell[    6334] = 32'h2f46587e;
    ram_cell[    6335] = 32'h477dac64;
    ram_cell[    6336] = 32'ha2df40b5;
    ram_cell[    6337] = 32'h7d3b2a1e;
    ram_cell[    6338] = 32'hd7c5ba7a;
    ram_cell[    6339] = 32'h25d81ead;
    ram_cell[    6340] = 32'heda44cea;
    ram_cell[    6341] = 32'h6ef60753;
    ram_cell[    6342] = 32'ha0d12bb9;
    ram_cell[    6343] = 32'h672bf5e1;
    ram_cell[    6344] = 32'h02d5562d;
    ram_cell[    6345] = 32'h913bc56c;
    ram_cell[    6346] = 32'hb159fb70;
    ram_cell[    6347] = 32'h52710028;
    ram_cell[    6348] = 32'h1b3d701a;
    ram_cell[    6349] = 32'h26f938a7;
    ram_cell[    6350] = 32'hc28e14db;
    ram_cell[    6351] = 32'ha54ab2ed;
    ram_cell[    6352] = 32'h430dceb6;
    ram_cell[    6353] = 32'hc7eedfe5;
    ram_cell[    6354] = 32'hb75e7912;
    ram_cell[    6355] = 32'h16889718;
    ram_cell[    6356] = 32'h60581294;
    ram_cell[    6357] = 32'h18277f8c;
    ram_cell[    6358] = 32'hfdedad97;
    ram_cell[    6359] = 32'h81b9172d;
    ram_cell[    6360] = 32'hc5d6bab7;
    ram_cell[    6361] = 32'h91d1d079;
    ram_cell[    6362] = 32'hadc5b366;
    ram_cell[    6363] = 32'h74f87c7e;
    ram_cell[    6364] = 32'h3a95125a;
    ram_cell[    6365] = 32'hc1284e4d;
    ram_cell[    6366] = 32'h766912ba;
    ram_cell[    6367] = 32'hb007d4fe;
    ram_cell[    6368] = 32'h4c3a1938;
    ram_cell[    6369] = 32'hdd05dbcc;
    ram_cell[    6370] = 32'he4985575;
    ram_cell[    6371] = 32'hf8fe8b14;
    ram_cell[    6372] = 32'h48b313c8;
    ram_cell[    6373] = 32'he85ad2e3;
    ram_cell[    6374] = 32'h5f0b574c;
    ram_cell[    6375] = 32'h9a986a0f;
    ram_cell[    6376] = 32'hfef1ee79;
    ram_cell[    6377] = 32'hbcf911f2;
    ram_cell[    6378] = 32'h7163845a;
    ram_cell[    6379] = 32'h3776bcd7;
    ram_cell[    6380] = 32'h9e91db4c;
    ram_cell[    6381] = 32'he99ff1df;
    ram_cell[    6382] = 32'he6c0e3ce;
    ram_cell[    6383] = 32'h4f90b2dc;
    ram_cell[    6384] = 32'h1050340d;
    ram_cell[    6385] = 32'h26310341;
    ram_cell[    6386] = 32'hf29c78a7;
    ram_cell[    6387] = 32'hde6d8a76;
    ram_cell[    6388] = 32'he0f2f9f7;
    ram_cell[    6389] = 32'h36e06f69;
    ram_cell[    6390] = 32'h92c110d4;
    ram_cell[    6391] = 32'hcc91ba22;
    ram_cell[    6392] = 32'he8eaa2a7;
    ram_cell[    6393] = 32'hbfe31d11;
    ram_cell[    6394] = 32'h6cfed26b;
    ram_cell[    6395] = 32'h17777f5f;
    ram_cell[    6396] = 32'hbeb2fee9;
    ram_cell[    6397] = 32'h47b5f3e1;
    ram_cell[    6398] = 32'hdee0aa6a;
    ram_cell[    6399] = 32'h4318a6a3;
    ram_cell[    6400] = 32'h80cbb6df;
    ram_cell[    6401] = 32'h28e504ae;
    ram_cell[    6402] = 32'h5f0e0d32;
    ram_cell[    6403] = 32'ha9673b77;
    ram_cell[    6404] = 32'hf4c7777c;
    ram_cell[    6405] = 32'hf1574f7f;
    ram_cell[    6406] = 32'h382637f5;
    ram_cell[    6407] = 32'h7feb966c;
    ram_cell[    6408] = 32'hd4b0518c;
    ram_cell[    6409] = 32'he6f161e2;
    ram_cell[    6410] = 32'h848ce970;
    ram_cell[    6411] = 32'hc9d52b7e;
    ram_cell[    6412] = 32'h98d4e717;
    ram_cell[    6413] = 32'he20f1bf6;
    ram_cell[    6414] = 32'h05f518ce;
    ram_cell[    6415] = 32'he0cba48b;
    ram_cell[    6416] = 32'hfafc076e;
    ram_cell[    6417] = 32'h9f666918;
    ram_cell[    6418] = 32'h02ee6209;
    ram_cell[    6419] = 32'h8eb90f7f;
    ram_cell[    6420] = 32'hed4e3d6b;
    ram_cell[    6421] = 32'h2920a804;
    ram_cell[    6422] = 32'hb463e484;
    ram_cell[    6423] = 32'ha06d9027;
    ram_cell[    6424] = 32'h2f2d6d37;
    ram_cell[    6425] = 32'h459f35b5;
    ram_cell[    6426] = 32'h0ad92b90;
    ram_cell[    6427] = 32'h20efdce2;
    ram_cell[    6428] = 32'hd1c9484b;
    ram_cell[    6429] = 32'h9e17dc89;
    ram_cell[    6430] = 32'hc569530c;
    ram_cell[    6431] = 32'h0b7df828;
    ram_cell[    6432] = 32'haaee6a86;
    ram_cell[    6433] = 32'he4c25228;
    ram_cell[    6434] = 32'h2b309279;
    ram_cell[    6435] = 32'h4b2d8a14;
    ram_cell[    6436] = 32'h0207523d;
    ram_cell[    6437] = 32'h3425d975;
    ram_cell[    6438] = 32'h16357467;
    ram_cell[    6439] = 32'h4ae2ed63;
    ram_cell[    6440] = 32'hb3ba39ac;
    ram_cell[    6441] = 32'ha2e63992;
    ram_cell[    6442] = 32'h391270fd;
    ram_cell[    6443] = 32'hca733f5f;
    ram_cell[    6444] = 32'haa24eb0f;
    ram_cell[    6445] = 32'h8daecf37;
    ram_cell[    6446] = 32'hba411e26;
    ram_cell[    6447] = 32'hc1ad89e1;
    ram_cell[    6448] = 32'h9707e93d;
    ram_cell[    6449] = 32'hea7b4b0d;
    ram_cell[    6450] = 32'hb6d4c16c;
    ram_cell[    6451] = 32'hf58279ae;
    ram_cell[    6452] = 32'hf7137c14;
    ram_cell[    6453] = 32'h85ba5331;
    ram_cell[    6454] = 32'hff41ac82;
    ram_cell[    6455] = 32'h4fab8b9e;
    ram_cell[    6456] = 32'he0e4568b;
    ram_cell[    6457] = 32'h698e569f;
    ram_cell[    6458] = 32'hdd34d895;
    ram_cell[    6459] = 32'hecf5de71;
    ram_cell[    6460] = 32'h9d019b21;
    ram_cell[    6461] = 32'h5945f0b9;
    ram_cell[    6462] = 32'h59748517;
    ram_cell[    6463] = 32'heb12b1f8;
    ram_cell[    6464] = 32'hd300a190;
    ram_cell[    6465] = 32'h7364f170;
    ram_cell[    6466] = 32'hbfa3eddf;
    ram_cell[    6467] = 32'h4269161a;
    ram_cell[    6468] = 32'hb6c01bfb;
    ram_cell[    6469] = 32'h7a7d1632;
    ram_cell[    6470] = 32'ha5b2d21b;
    ram_cell[    6471] = 32'head28657;
    ram_cell[    6472] = 32'h8b083cd8;
    ram_cell[    6473] = 32'h5f30295b;
    ram_cell[    6474] = 32'h679b675a;
    ram_cell[    6475] = 32'h5c140a75;
    ram_cell[    6476] = 32'hfb836c1e;
    ram_cell[    6477] = 32'h2dc49c52;
    ram_cell[    6478] = 32'hf8b7cb52;
    ram_cell[    6479] = 32'h1366e676;
    ram_cell[    6480] = 32'h96e19491;
    ram_cell[    6481] = 32'h115474ac;
    ram_cell[    6482] = 32'hb4fdb76a;
    ram_cell[    6483] = 32'he830f8a5;
    ram_cell[    6484] = 32'h88e85787;
    ram_cell[    6485] = 32'h980b5e3c;
    ram_cell[    6486] = 32'hd4ce4b0d;
    ram_cell[    6487] = 32'hee89b7d0;
    ram_cell[    6488] = 32'h699e927b;
    ram_cell[    6489] = 32'he3e3e75a;
    ram_cell[    6490] = 32'ha356bf97;
    ram_cell[    6491] = 32'h2568916f;
    ram_cell[    6492] = 32'h78accb67;
    ram_cell[    6493] = 32'h04b6ffb9;
    ram_cell[    6494] = 32'h82d7170f;
    ram_cell[    6495] = 32'h78252dad;
    ram_cell[    6496] = 32'h53340f38;
    ram_cell[    6497] = 32'h7d502e15;
    ram_cell[    6498] = 32'h9494edd8;
    ram_cell[    6499] = 32'hd2a20763;
    ram_cell[    6500] = 32'h6148bc53;
    ram_cell[    6501] = 32'hf142c55e;
    ram_cell[    6502] = 32'h21861f52;
    ram_cell[    6503] = 32'h5ce31b2d;
    ram_cell[    6504] = 32'hb170abf8;
    ram_cell[    6505] = 32'h1c0c0fa0;
    ram_cell[    6506] = 32'hba533167;
    ram_cell[    6507] = 32'h6cc419b9;
    ram_cell[    6508] = 32'hc44079f6;
    ram_cell[    6509] = 32'h7917aa42;
    ram_cell[    6510] = 32'h9db8029e;
    ram_cell[    6511] = 32'hc019393f;
    ram_cell[    6512] = 32'h26bdc761;
    ram_cell[    6513] = 32'h0c2ae080;
    ram_cell[    6514] = 32'h152a7212;
    ram_cell[    6515] = 32'ha0f508f8;
    ram_cell[    6516] = 32'h596cd463;
    ram_cell[    6517] = 32'h9c236137;
    ram_cell[    6518] = 32'hf97c93be;
    ram_cell[    6519] = 32'h573aedb0;
    ram_cell[    6520] = 32'hbca7ea8f;
    ram_cell[    6521] = 32'h35b3f9da;
    ram_cell[    6522] = 32'ha39c685a;
    ram_cell[    6523] = 32'h3c7fc846;
    ram_cell[    6524] = 32'ha1177122;
    ram_cell[    6525] = 32'h04f36567;
    ram_cell[    6526] = 32'h5236af22;
    ram_cell[    6527] = 32'h3cd3ab01;
    ram_cell[    6528] = 32'h5410f7a7;
    ram_cell[    6529] = 32'h67c62783;
    ram_cell[    6530] = 32'hddc09e76;
    ram_cell[    6531] = 32'h66770bc7;
    ram_cell[    6532] = 32'hc2bbf2ea;
    ram_cell[    6533] = 32'h4161327c;
    ram_cell[    6534] = 32'h6c809fbe;
    ram_cell[    6535] = 32'h1561c768;
    ram_cell[    6536] = 32'h71d4afe3;
    ram_cell[    6537] = 32'h5b237c71;
    ram_cell[    6538] = 32'h95bf6339;
    ram_cell[    6539] = 32'h4856dcf0;
    ram_cell[    6540] = 32'h128ca186;
    ram_cell[    6541] = 32'hebaf1639;
    ram_cell[    6542] = 32'h27b80347;
    ram_cell[    6543] = 32'h45d3fc6a;
    ram_cell[    6544] = 32'hc9b99120;
    ram_cell[    6545] = 32'hc1becbf0;
    ram_cell[    6546] = 32'hd69fffa3;
    ram_cell[    6547] = 32'had20eec7;
    ram_cell[    6548] = 32'hc1957b95;
    ram_cell[    6549] = 32'hd0d7e56b;
    ram_cell[    6550] = 32'h2d03f4dd;
    ram_cell[    6551] = 32'h16a947d2;
    ram_cell[    6552] = 32'hca1cb944;
    ram_cell[    6553] = 32'h824fc5fa;
    ram_cell[    6554] = 32'hbdc18376;
    ram_cell[    6555] = 32'habd0fe18;
    ram_cell[    6556] = 32'h40767259;
    ram_cell[    6557] = 32'h42465184;
    ram_cell[    6558] = 32'h2662e92a;
    ram_cell[    6559] = 32'hc86fbbeb;
    ram_cell[    6560] = 32'hc0e6d975;
    ram_cell[    6561] = 32'h5ab1e038;
    ram_cell[    6562] = 32'h349c01b2;
    ram_cell[    6563] = 32'he3a03468;
    ram_cell[    6564] = 32'h0867a054;
    ram_cell[    6565] = 32'hda2cfff6;
    ram_cell[    6566] = 32'h073b7233;
    ram_cell[    6567] = 32'h5fabaea2;
    ram_cell[    6568] = 32'h51038131;
    ram_cell[    6569] = 32'h7d62f212;
    ram_cell[    6570] = 32'h288930dc;
    ram_cell[    6571] = 32'hc01e9d90;
    ram_cell[    6572] = 32'h7bf8e47e;
    ram_cell[    6573] = 32'hc422a54a;
    ram_cell[    6574] = 32'h7d0a7935;
    ram_cell[    6575] = 32'h7155e87f;
    ram_cell[    6576] = 32'h1e2a25e2;
    ram_cell[    6577] = 32'hf8a3abca;
    ram_cell[    6578] = 32'hd6bcf684;
    ram_cell[    6579] = 32'h2b84810b;
    ram_cell[    6580] = 32'h24fc693e;
    ram_cell[    6581] = 32'h2f7c59e3;
    ram_cell[    6582] = 32'h7181d2ae;
    ram_cell[    6583] = 32'hcd751063;
    ram_cell[    6584] = 32'hcc1282df;
    ram_cell[    6585] = 32'h7beb52e4;
    ram_cell[    6586] = 32'h16638930;
    ram_cell[    6587] = 32'h8f0787c0;
    ram_cell[    6588] = 32'hd840e11f;
    ram_cell[    6589] = 32'h7771ee28;
    ram_cell[    6590] = 32'h4d56df8a;
    ram_cell[    6591] = 32'h9ad3b623;
    ram_cell[    6592] = 32'h27f4873d;
    ram_cell[    6593] = 32'h03934c3a;
    ram_cell[    6594] = 32'ha3ce52a0;
    ram_cell[    6595] = 32'h3db1aea3;
    ram_cell[    6596] = 32'h1dc79805;
    ram_cell[    6597] = 32'hb2978a13;
    ram_cell[    6598] = 32'h0685cde1;
    ram_cell[    6599] = 32'hee0e414d;
    ram_cell[    6600] = 32'h3475f76a;
    ram_cell[    6601] = 32'h90db71bd;
    ram_cell[    6602] = 32'hfdda57af;
    ram_cell[    6603] = 32'hb96cdf0f;
    ram_cell[    6604] = 32'ha760c341;
    ram_cell[    6605] = 32'h4858ed0c;
    ram_cell[    6606] = 32'h7f5de164;
    ram_cell[    6607] = 32'h8f32da7e;
    ram_cell[    6608] = 32'h9a2d470d;
    ram_cell[    6609] = 32'hd48a33d1;
    ram_cell[    6610] = 32'h117e00f5;
    ram_cell[    6611] = 32'h4bf05904;
    ram_cell[    6612] = 32'h906966b5;
    ram_cell[    6613] = 32'hec34192a;
    ram_cell[    6614] = 32'h73b6ffe3;
    ram_cell[    6615] = 32'hd2290119;
    ram_cell[    6616] = 32'h72511a4b;
    ram_cell[    6617] = 32'h7489c56e;
    ram_cell[    6618] = 32'h247b4183;
    ram_cell[    6619] = 32'h8b5f9218;
    ram_cell[    6620] = 32'h90896873;
    ram_cell[    6621] = 32'hbeb2b146;
    ram_cell[    6622] = 32'h7dc61fe4;
    ram_cell[    6623] = 32'h827772da;
    ram_cell[    6624] = 32'h906dd728;
    ram_cell[    6625] = 32'h2b6cf20d;
    ram_cell[    6626] = 32'h44f5993a;
    ram_cell[    6627] = 32'h9aa3181d;
    ram_cell[    6628] = 32'h606a471c;
    ram_cell[    6629] = 32'h61151835;
    ram_cell[    6630] = 32'hc23ba287;
    ram_cell[    6631] = 32'h6417df1e;
    ram_cell[    6632] = 32'h7c080228;
    ram_cell[    6633] = 32'hc42cc800;
    ram_cell[    6634] = 32'h4443d016;
    ram_cell[    6635] = 32'h270885e7;
    ram_cell[    6636] = 32'he411fc55;
    ram_cell[    6637] = 32'ha1203525;
    ram_cell[    6638] = 32'h9fa834cb;
    ram_cell[    6639] = 32'h3f0e0a01;
    ram_cell[    6640] = 32'hd0f9ab77;
    ram_cell[    6641] = 32'h5f9cbbc4;
    ram_cell[    6642] = 32'h8da12892;
    ram_cell[    6643] = 32'hd21cc7dd;
    ram_cell[    6644] = 32'h8e6fdaee;
    ram_cell[    6645] = 32'hc9bb6767;
    ram_cell[    6646] = 32'h6ee88168;
    ram_cell[    6647] = 32'hd3cde972;
    ram_cell[    6648] = 32'h6e1443d2;
    ram_cell[    6649] = 32'h513f44e1;
    ram_cell[    6650] = 32'h7303881c;
    ram_cell[    6651] = 32'h15ae1886;
    ram_cell[    6652] = 32'h061576ee;
    ram_cell[    6653] = 32'h0cffe473;
    ram_cell[    6654] = 32'h9ba92663;
    ram_cell[    6655] = 32'h07aa184a;
    ram_cell[    6656] = 32'h4936a603;
    ram_cell[    6657] = 32'h6e62ccc9;
    ram_cell[    6658] = 32'ha9ff3da0;
    ram_cell[    6659] = 32'hc42f47de;
    ram_cell[    6660] = 32'ha9b60f11;
    ram_cell[    6661] = 32'hf631344d;
    ram_cell[    6662] = 32'hc98d36ff;
    ram_cell[    6663] = 32'h444415cb;
    ram_cell[    6664] = 32'h396543fd;
    ram_cell[    6665] = 32'h0cdc2620;
    ram_cell[    6666] = 32'ha20bae14;
    ram_cell[    6667] = 32'hb99176ae;
    ram_cell[    6668] = 32'hee6c1ab8;
    ram_cell[    6669] = 32'h5397bd6e;
    ram_cell[    6670] = 32'h1bff0dc3;
    ram_cell[    6671] = 32'hb97e9d49;
    ram_cell[    6672] = 32'h107eca42;
    ram_cell[    6673] = 32'h7b5c9515;
    ram_cell[    6674] = 32'hfd7a78ea;
    ram_cell[    6675] = 32'h3bef0ac2;
    ram_cell[    6676] = 32'h3fa35512;
    ram_cell[    6677] = 32'h2205449c;
    ram_cell[    6678] = 32'haf02fca6;
    ram_cell[    6679] = 32'hb951fece;
    ram_cell[    6680] = 32'h99511e49;
    ram_cell[    6681] = 32'hbc614cd8;
    ram_cell[    6682] = 32'h22308d0f;
    ram_cell[    6683] = 32'hc597cc0f;
    ram_cell[    6684] = 32'h338f5a2c;
    ram_cell[    6685] = 32'hb253f324;
    ram_cell[    6686] = 32'ha6963ca2;
    ram_cell[    6687] = 32'h120f098c;
    ram_cell[    6688] = 32'ha350fc89;
    ram_cell[    6689] = 32'h9f69d8b3;
    ram_cell[    6690] = 32'h375d28ac;
    ram_cell[    6691] = 32'h207fe172;
    ram_cell[    6692] = 32'h59ce8205;
    ram_cell[    6693] = 32'h779f80ca;
    ram_cell[    6694] = 32'h9dd7a83a;
    ram_cell[    6695] = 32'hfb172aa7;
    ram_cell[    6696] = 32'h150f2c94;
    ram_cell[    6697] = 32'h85fdf711;
    ram_cell[    6698] = 32'h4b7deb1d;
    ram_cell[    6699] = 32'h89aa5120;
    ram_cell[    6700] = 32'hb4d47cf2;
    ram_cell[    6701] = 32'h61004bc0;
    ram_cell[    6702] = 32'hfd6f61bd;
    ram_cell[    6703] = 32'ha3dd36d3;
    ram_cell[    6704] = 32'h5b95591a;
    ram_cell[    6705] = 32'h685e3607;
    ram_cell[    6706] = 32'h0f9aa920;
    ram_cell[    6707] = 32'he4e0c8af;
    ram_cell[    6708] = 32'h80af95fe;
    ram_cell[    6709] = 32'h11ef057a;
    ram_cell[    6710] = 32'h9cf2780f;
    ram_cell[    6711] = 32'h161f03f5;
    ram_cell[    6712] = 32'h178df102;
    ram_cell[    6713] = 32'h96da5de9;
    ram_cell[    6714] = 32'h1a469292;
    ram_cell[    6715] = 32'h02d708e2;
    ram_cell[    6716] = 32'h1465328b;
    ram_cell[    6717] = 32'h63d53ce2;
    ram_cell[    6718] = 32'hd26672a5;
    ram_cell[    6719] = 32'h6453ec76;
    ram_cell[    6720] = 32'h7cefe2db;
    ram_cell[    6721] = 32'h03a6030b;
    ram_cell[    6722] = 32'h43236b78;
    ram_cell[    6723] = 32'h7dbb20f6;
    ram_cell[    6724] = 32'h174dd518;
    ram_cell[    6725] = 32'haeaca10c;
    ram_cell[    6726] = 32'haef0950a;
    ram_cell[    6727] = 32'h7e6f8ba7;
    ram_cell[    6728] = 32'hfb2e24a5;
    ram_cell[    6729] = 32'h240f3973;
    ram_cell[    6730] = 32'h4eca69f4;
    ram_cell[    6731] = 32'h829010b6;
    ram_cell[    6732] = 32'h035d41c8;
    ram_cell[    6733] = 32'hd2d463eb;
    ram_cell[    6734] = 32'he51dddce;
    ram_cell[    6735] = 32'hb75a2015;
    ram_cell[    6736] = 32'hd948fa65;
    ram_cell[    6737] = 32'hcbec5fc1;
    ram_cell[    6738] = 32'ha6391d6d;
    ram_cell[    6739] = 32'hb2728cb5;
    ram_cell[    6740] = 32'h09f19f2b;
    ram_cell[    6741] = 32'hf9f2d47d;
    ram_cell[    6742] = 32'h7bfac8fd;
    ram_cell[    6743] = 32'hcd461167;
    ram_cell[    6744] = 32'h7a77a920;
    ram_cell[    6745] = 32'h57141db7;
    ram_cell[    6746] = 32'ha317b7aa;
    ram_cell[    6747] = 32'h9e52f67d;
    ram_cell[    6748] = 32'hfdf445d5;
    ram_cell[    6749] = 32'hd05d0bc8;
    ram_cell[    6750] = 32'ha3c5bc3d;
    ram_cell[    6751] = 32'h7b22d95c;
    ram_cell[    6752] = 32'hf781fb96;
    ram_cell[    6753] = 32'heb4232e3;
    ram_cell[    6754] = 32'h3b753c6a;
    ram_cell[    6755] = 32'hd292df30;
    ram_cell[    6756] = 32'h02cfa32e;
    ram_cell[    6757] = 32'h00e5107b;
    ram_cell[    6758] = 32'hf3781429;
    ram_cell[    6759] = 32'h814f0608;
    ram_cell[    6760] = 32'h84210d5c;
    ram_cell[    6761] = 32'h57093bf9;
    ram_cell[    6762] = 32'h6f7a8a1b;
    ram_cell[    6763] = 32'h4071ad1a;
    ram_cell[    6764] = 32'ha3d4a8ec;
    ram_cell[    6765] = 32'hc886efcd;
    ram_cell[    6766] = 32'h075e1fa5;
    ram_cell[    6767] = 32'h922f0692;
    ram_cell[    6768] = 32'hd51f2550;
    ram_cell[    6769] = 32'he5f3d6d8;
    ram_cell[    6770] = 32'hadae50a0;
    ram_cell[    6771] = 32'h3246ba07;
    ram_cell[    6772] = 32'h10103263;
    ram_cell[    6773] = 32'h3161d03c;
    ram_cell[    6774] = 32'hcbaca96b;
    ram_cell[    6775] = 32'hb38a2caf;
    ram_cell[    6776] = 32'h39452dab;
    ram_cell[    6777] = 32'h0b00a775;
    ram_cell[    6778] = 32'h8e03c596;
    ram_cell[    6779] = 32'h4df72566;
    ram_cell[    6780] = 32'h44b23beb;
    ram_cell[    6781] = 32'h520ac382;
    ram_cell[    6782] = 32'h4ec5c871;
    ram_cell[    6783] = 32'he0a64c40;
    ram_cell[    6784] = 32'h9adb0710;
    ram_cell[    6785] = 32'h495b184d;
    ram_cell[    6786] = 32'h28294b76;
    ram_cell[    6787] = 32'hfa7c360a;
    ram_cell[    6788] = 32'h38e25d80;
    ram_cell[    6789] = 32'hcd2ba1a4;
    ram_cell[    6790] = 32'h72372edb;
    ram_cell[    6791] = 32'hea6f9279;
    ram_cell[    6792] = 32'h26f6a82d;
    ram_cell[    6793] = 32'h89a4bdc0;
    ram_cell[    6794] = 32'hf1a2d15f;
    ram_cell[    6795] = 32'h287f91c9;
    ram_cell[    6796] = 32'h491c0d1e;
    ram_cell[    6797] = 32'h8a5e7eae;
    ram_cell[    6798] = 32'ha643dabb;
    ram_cell[    6799] = 32'h2c1669c1;
    ram_cell[    6800] = 32'hf36e9ac3;
    ram_cell[    6801] = 32'h0bb951fb;
    ram_cell[    6802] = 32'h1b8eec4b;
    ram_cell[    6803] = 32'hba2a85f5;
    ram_cell[    6804] = 32'hb6e3008d;
    ram_cell[    6805] = 32'h6391dd08;
    ram_cell[    6806] = 32'h598a71f6;
    ram_cell[    6807] = 32'h1118f70e;
    ram_cell[    6808] = 32'hb4e22dfa;
    ram_cell[    6809] = 32'hb548522c;
    ram_cell[    6810] = 32'hb504d66a;
    ram_cell[    6811] = 32'h5fb7fe04;
    ram_cell[    6812] = 32'hae93bd7b;
    ram_cell[    6813] = 32'hf45a5453;
    ram_cell[    6814] = 32'h986814c0;
    ram_cell[    6815] = 32'hdf4690e8;
    ram_cell[    6816] = 32'hc15cae1a;
    ram_cell[    6817] = 32'h598b11a2;
    ram_cell[    6818] = 32'h26e078bf;
    ram_cell[    6819] = 32'hdea7ee5c;
    ram_cell[    6820] = 32'h0768a027;
    ram_cell[    6821] = 32'h2dc65c4a;
    ram_cell[    6822] = 32'h623536bc;
    ram_cell[    6823] = 32'h242f7a7a;
    ram_cell[    6824] = 32'hc367887c;
    ram_cell[    6825] = 32'h1df88bd7;
    ram_cell[    6826] = 32'hc3e5db2f;
    ram_cell[    6827] = 32'hd25864cd;
    ram_cell[    6828] = 32'h5409446f;
    ram_cell[    6829] = 32'hfb0e86a4;
    ram_cell[    6830] = 32'h01f52609;
    ram_cell[    6831] = 32'h83bdd81f;
    ram_cell[    6832] = 32'ha7217cc8;
    ram_cell[    6833] = 32'hafe5a8d8;
    ram_cell[    6834] = 32'h2e4a36a2;
    ram_cell[    6835] = 32'h56309b12;
    ram_cell[    6836] = 32'hf3869ec1;
    ram_cell[    6837] = 32'h01711ab1;
    ram_cell[    6838] = 32'h992dc4ec;
    ram_cell[    6839] = 32'h4b31fd65;
    ram_cell[    6840] = 32'he93033f5;
    ram_cell[    6841] = 32'hd46162cf;
    ram_cell[    6842] = 32'he1fffe88;
    ram_cell[    6843] = 32'hb36fcc7e;
    ram_cell[    6844] = 32'hdda52766;
    ram_cell[    6845] = 32'h44775257;
    ram_cell[    6846] = 32'h287d98f9;
    ram_cell[    6847] = 32'h3b93bb21;
    ram_cell[    6848] = 32'hda356dc5;
    ram_cell[    6849] = 32'h86bfe4c2;
    ram_cell[    6850] = 32'h605fc284;
    ram_cell[    6851] = 32'h28543de7;
    ram_cell[    6852] = 32'h77de41e0;
    ram_cell[    6853] = 32'h5e9c3857;
    ram_cell[    6854] = 32'hf9f2b989;
    ram_cell[    6855] = 32'hd6cbe50d;
    ram_cell[    6856] = 32'hd8b88ea0;
    ram_cell[    6857] = 32'hacba00df;
    ram_cell[    6858] = 32'h2f90671d;
    ram_cell[    6859] = 32'hb6bb5370;
    ram_cell[    6860] = 32'h13ae75bc;
    ram_cell[    6861] = 32'hb95c2ef7;
    ram_cell[    6862] = 32'h4c2ebbd7;
    ram_cell[    6863] = 32'hb9228872;
    ram_cell[    6864] = 32'h122b9410;
    ram_cell[    6865] = 32'hf1efa8b4;
    ram_cell[    6866] = 32'h1ee100ac;
    ram_cell[    6867] = 32'h07145dd7;
    ram_cell[    6868] = 32'hcf74689c;
    ram_cell[    6869] = 32'h9039e6c0;
    ram_cell[    6870] = 32'h89cee294;
    ram_cell[    6871] = 32'h7c9e7235;
    ram_cell[    6872] = 32'ha1a01709;
    ram_cell[    6873] = 32'hb30cb819;
    ram_cell[    6874] = 32'hf5bf226d;
    ram_cell[    6875] = 32'hc44f4289;
    ram_cell[    6876] = 32'h8741c78c;
    ram_cell[    6877] = 32'h82759f2f;
    ram_cell[    6878] = 32'h1a2bc94b;
    ram_cell[    6879] = 32'h119cab1e;
    ram_cell[    6880] = 32'h3aa61102;
    ram_cell[    6881] = 32'hce775099;
    ram_cell[    6882] = 32'hf188d344;
    ram_cell[    6883] = 32'hf653a3e6;
    ram_cell[    6884] = 32'h7c512b7d;
    ram_cell[    6885] = 32'hee93c924;
    ram_cell[    6886] = 32'he929b6bc;
    ram_cell[    6887] = 32'h6fc541aa;
    ram_cell[    6888] = 32'hfb16ebe2;
    ram_cell[    6889] = 32'hc829137a;
    ram_cell[    6890] = 32'h1c19a839;
    ram_cell[    6891] = 32'h0b179869;
    ram_cell[    6892] = 32'h15e19bbc;
    ram_cell[    6893] = 32'hbf1ab06b;
    ram_cell[    6894] = 32'h6ff869f7;
    ram_cell[    6895] = 32'hd3edb561;
    ram_cell[    6896] = 32'hb25d3e3f;
    ram_cell[    6897] = 32'hf4e65ee8;
    ram_cell[    6898] = 32'h26fe5ec1;
    ram_cell[    6899] = 32'ha4a54ee1;
    ram_cell[    6900] = 32'h14c711f8;
    ram_cell[    6901] = 32'ha6d54f21;
    ram_cell[    6902] = 32'h6f60a43d;
    ram_cell[    6903] = 32'hf257e838;
    ram_cell[    6904] = 32'h6738488e;
    ram_cell[    6905] = 32'h0c7cda43;
    ram_cell[    6906] = 32'hb643b4de;
    ram_cell[    6907] = 32'heb3b6e3f;
    ram_cell[    6908] = 32'h9e232312;
    ram_cell[    6909] = 32'hed6dbf29;
    ram_cell[    6910] = 32'h713ffe03;
    ram_cell[    6911] = 32'h004dea6e;
    ram_cell[    6912] = 32'he3fd81e1;
    ram_cell[    6913] = 32'hed2a2c8f;
    ram_cell[    6914] = 32'h7e5f0050;
    ram_cell[    6915] = 32'h598900cd;
    ram_cell[    6916] = 32'hb2934b1e;
    ram_cell[    6917] = 32'h04f9d5ca;
    ram_cell[    6918] = 32'h08cff6e2;
    ram_cell[    6919] = 32'h9495b6a3;
    ram_cell[    6920] = 32'h27d82fec;
    ram_cell[    6921] = 32'h1291a98a;
    ram_cell[    6922] = 32'h66a6d80b;
    ram_cell[    6923] = 32'haf4eef01;
    ram_cell[    6924] = 32'hf6198f7a;
    ram_cell[    6925] = 32'h59bfa876;
    ram_cell[    6926] = 32'h561c1dd8;
    ram_cell[    6927] = 32'h355a87fd;
    ram_cell[    6928] = 32'hf5680f12;
    ram_cell[    6929] = 32'hd65a71e3;
    ram_cell[    6930] = 32'h8c62c33e;
    ram_cell[    6931] = 32'h4f53833c;
    ram_cell[    6932] = 32'h1a2c041d;
    ram_cell[    6933] = 32'h6c1ae18a;
    ram_cell[    6934] = 32'h72fdf358;
    ram_cell[    6935] = 32'hd7b6e8f3;
    ram_cell[    6936] = 32'hf3ca2dae;
    ram_cell[    6937] = 32'h08d14ad4;
    ram_cell[    6938] = 32'had3db350;
    ram_cell[    6939] = 32'hebdfa976;
    ram_cell[    6940] = 32'h8a2d2baf;
    ram_cell[    6941] = 32'hc185459e;
    ram_cell[    6942] = 32'h92ae8a3a;
    ram_cell[    6943] = 32'hf64709d3;
    ram_cell[    6944] = 32'h4f1c1654;
    ram_cell[    6945] = 32'h5d28892e;
    ram_cell[    6946] = 32'hf5061739;
    ram_cell[    6947] = 32'hf8e51e0b;
    ram_cell[    6948] = 32'haf8f88ad;
    ram_cell[    6949] = 32'h3c1e5083;
    ram_cell[    6950] = 32'h2af097d3;
    ram_cell[    6951] = 32'h2a0c474f;
    ram_cell[    6952] = 32'hfc955b37;
    ram_cell[    6953] = 32'h055e70c9;
    ram_cell[    6954] = 32'hd70765fb;
    ram_cell[    6955] = 32'hb07ffff0;
    ram_cell[    6956] = 32'h19a71cd5;
    ram_cell[    6957] = 32'h0deb0ae3;
    ram_cell[    6958] = 32'he4a6b36c;
    ram_cell[    6959] = 32'hb15033a7;
    ram_cell[    6960] = 32'haea39a4a;
    ram_cell[    6961] = 32'h06982b33;
    ram_cell[    6962] = 32'hf5c982ff;
    ram_cell[    6963] = 32'h1f820d39;
    ram_cell[    6964] = 32'h61842951;
    ram_cell[    6965] = 32'hbac0ca4e;
    ram_cell[    6966] = 32'h7dc3afa4;
    ram_cell[    6967] = 32'hef450c55;
    ram_cell[    6968] = 32'h8cc4de6c;
    ram_cell[    6969] = 32'h59ff387a;
    ram_cell[    6970] = 32'h63a6f9ea;
    ram_cell[    6971] = 32'h9b06a254;
    ram_cell[    6972] = 32'h8b12d1cf;
    ram_cell[    6973] = 32'hc5834ff3;
    ram_cell[    6974] = 32'hf4992e15;
    ram_cell[    6975] = 32'h8891a9e7;
    ram_cell[    6976] = 32'h2ad8cd96;
    ram_cell[    6977] = 32'hd28fa600;
    ram_cell[    6978] = 32'hd1c43ec8;
    ram_cell[    6979] = 32'hcd4d9a79;
    ram_cell[    6980] = 32'hbc4a4cf3;
    ram_cell[    6981] = 32'ha8a80c47;
    ram_cell[    6982] = 32'hdff552f2;
    ram_cell[    6983] = 32'h52b20425;
    ram_cell[    6984] = 32'h1b8e7227;
    ram_cell[    6985] = 32'h8b8ca22e;
    ram_cell[    6986] = 32'he34cce54;
    ram_cell[    6987] = 32'h9977ba2f;
    ram_cell[    6988] = 32'h14c69e6a;
    ram_cell[    6989] = 32'h66c0f5f3;
    ram_cell[    6990] = 32'h6a25537c;
    ram_cell[    6991] = 32'he57747d2;
    ram_cell[    6992] = 32'h226eedb4;
    ram_cell[    6993] = 32'hb517b538;
    ram_cell[    6994] = 32'hdf3e861b;
    ram_cell[    6995] = 32'ha8497fb7;
    ram_cell[    6996] = 32'he2971565;
    ram_cell[    6997] = 32'haa0afb11;
    ram_cell[    6998] = 32'h564192b4;
    ram_cell[    6999] = 32'hf1563f80;
    ram_cell[    7000] = 32'hd1b58ca4;
    ram_cell[    7001] = 32'hb1e8e5bd;
    ram_cell[    7002] = 32'h2551a9bb;
    ram_cell[    7003] = 32'h4db29f2a;
    ram_cell[    7004] = 32'h7d261d92;
    ram_cell[    7005] = 32'h5b571d14;
    ram_cell[    7006] = 32'hbdcfae6c;
    ram_cell[    7007] = 32'h46a147bc;
    ram_cell[    7008] = 32'h8a6c26b2;
    ram_cell[    7009] = 32'ha51512e4;
    ram_cell[    7010] = 32'h947568ad;
    ram_cell[    7011] = 32'hbc17e687;
    ram_cell[    7012] = 32'h162296d2;
    ram_cell[    7013] = 32'he3ffd384;
    ram_cell[    7014] = 32'h3b0aa58f;
    ram_cell[    7015] = 32'hc6871b74;
    ram_cell[    7016] = 32'hf8e4e510;
    ram_cell[    7017] = 32'h50b84614;
    ram_cell[    7018] = 32'hb63aa539;
    ram_cell[    7019] = 32'h7872fcb3;
    ram_cell[    7020] = 32'h940677ed;
    ram_cell[    7021] = 32'ha5ec66b0;
    ram_cell[    7022] = 32'h52bc6b6c;
    ram_cell[    7023] = 32'hbcf6cc94;
    ram_cell[    7024] = 32'heb66c070;
    ram_cell[    7025] = 32'h52f17991;
    ram_cell[    7026] = 32'hf4911ef7;
    ram_cell[    7027] = 32'haec89288;
    ram_cell[    7028] = 32'hcc3c4ecb;
    ram_cell[    7029] = 32'hfd1d08c3;
    ram_cell[    7030] = 32'hb8285339;
    ram_cell[    7031] = 32'h423401e9;
    ram_cell[    7032] = 32'h095030c6;
    ram_cell[    7033] = 32'h0542586c;
    ram_cell[    7034] = 32'h462ff673;
    ram_cell[    7035] = 32'h634ba7a7;
    ram_cell[    7036] = 32'h98dfb682;
    ram_cell[    7037] = 32'hd029d6db;
    ram_cell[    7038] = 32'h7bc1c9a4;
    ram_cell[    7039] = 32'hc73931a1;
    ram_cell[    7040] = 32'hd9714bfa;
    ram_cell[    7041] = 32'ha37bebc1;
    ram_cell[    7042] = 32'hc38dfaf3;
    ram_cell[    7043] = 32'h1e27e3ee;
    ram_cell[    7044] = 32'h7182d2f9;
    ram_cell[    7045] = 32'hcbfa55da;
    ram_cell[    7046] = 32'ha094644e;
    ram_cell[    7047] = 32'hf58f211e;
    ram_cell[    7048] = 32'haa1ccfb2;
    ram_cell[    7049] = 32'hbccc9992;
    ram_cell[    7050] = 32'hc244ef23;
    ram_cell[    7051] = 32'h2b814fa2;
    ram_cell[    7052] = 32'hfab0e7b0;
    ram_cell[    7053] = 32'h3c8c31a5;
    ram_cell[    7054] = 32'hec166e4c;
    ram_cell[    7055] = 32'h9e9ed0b7;
    ram_cell[    7056] = 32'h5053f821;
    ram_cell[    7057] = 32'he1b5adcc;
    ram_cell[    7058] = 32'hc8d48ccf;
    ram_cell[    7059] = 32'h99c47255;
    ram_cell[    7060] = 32'h34944dfe;
    ram_cell[    7061] = 32'ha3639f4b;
    ram_cell[    7062] = 32'hf3cf3b03;
    ram_cell[    7063] = 32'he6ae157f;
    ram_cell[    7064] = 32'heabdd4de;
    ram_cell[    7065] = 32'h7bd5212e;
    ram_cell[    7066] = 32'hfdda771e;
    ram_cell[    7067] = 32'h5aacd810;
    ram_cell[    7068] = 32'h7090615c;
    ram_cell[    7069] = 32'hb0d9b2ae;
    ram_cell[    7070] = 32'hd61a7d42;
    ram_cell[    7071] = 32'hd1ca0eef;
    ram_cell[    7072] = 32'h65e42d6a;
    ram_cell[    7073] = 32'hc01177df;
    ram_cell[    7074] = 32'h2dfa8c2b;
    ram_cell[    7075] = 32'hf8e2fadd;
    ram_cell[    7076] = 32'h84623698;
    ram_cell[    7077] = 32'hb1d2282f;
    ram_cell[    7078] = 32'h44944bd2;
    ram_cell[    7079] = 32'h04227ac8;
    ram_cell[    7080] = 32'he3b6e65f;
    ram_cell[    7081] = 32'h89b3c4a2;
    ram_cell[    7082] = 32'h9ffc4ff9;
    ram_cell[    7083] = 32'hfe3ee5dc;
    ram_cell[    7084] = 32'hd3893df8;
    ram_cell[    7085] = 32'hf601ef68;
    ram_cell[    7086] = 32'h769b9fa7;
    ram_cell[    7087] = 32'hd6f06c71;
    ram_cell[    7088] = 32'hff0369ac;
    ram_cell[    7089] = 32'h3bf1dbd8;
    ram_cell[    7090] = 32'h31096c5d;
    ram_cell[    7091] = 32'hd9fcdbac;
    ram_cell[    7092] = 32'h53787d1b;
    ram_cell[    7093] = 32'hd99527b6;
    ram_cell[    7094] = 32'hd2ce797e;
    ram_cell[    7095] = 32'hae70ff0e;
    ram_cell[    7096] = 32'h92b1e5b5;
    ram_cell[    7097] = 32'h13436137;
    ram_cell[    7098] = 32'h362811f8;
    ram_cell[    7099] = 32'h52bd5523;
    ram_cell[    7100] = 32'h30cea4f1;
    ram_cell[    7101] = 32'hfa400ecf;
    ram_cell[    7102] = 32'h526d1be7;
    ram_cell[    7103] = 32'hf6f25101;
    ram_cell[    7104] = 32'hf40f47bd;
    ram_cell[    7105] = 32'h5b273d4d;
    ram_cell[    7106] = 32'h06a82948;
    ram_cell[    7107] = 32'h9ef79fa7;
    ram_cell[    7108] = 32'hc9f3f609;
    ram_cell[    7109] = 32'hed606e86;
    ram_cell[    7110] = 32'h6f7f00b0;
    ram_cell[    7111] = 32'hcc9f7b01;
    ram_cell[    7112] = 32'hef5c9e9f;
    ram_cell[    7113] = 32'h9fe71baf;
    ram_cell[    7114] = 32'hf16ec73b;
    ram_cell[    7115] = 32'hd08ece95;
    ram_cell[    7116] = 32'hd39268af;
    ram_cell[    7117] = 32'h3ebc8d0c;
    ram_cell[    7118] = 32'h92ead91b;
    ram_cell[    7119] = 32'h64b6632a;
    ram_cell[    7120] = 32'h57e4a45e;
    ram_cell[    7121] = 32'hd7a6fd2d;
    ram_cell[    7122] = 32'h84b1f736;
    ram_cell[    7123] = 32'h7deea4f8;
    ram_cell[    7124] = 32'he04e2b0e;
    ram_cell[    7125] = 32'hd27eb091;
    ram_cell[    7126] = 32'h1e4df0ef;
    ram_cell[    7127] = 32'h8ad6a3fd;
    ram_cell[    7128] = 32'h4a8f0842;
    ram_cell[    7129] = 32'h0e8aa592;
    ram_cell[    7130] = 32'h9d22270e;
    ram_cell[    7131] = 32'h8a42ea6b;
    ram_cell[    7132] = 32'hcdc2d0b3;
    ram_cell[    7133] = 32'h8d03aa89;
    ram_cell[    7134] = 32'hd4d37ae8;
    ram_cell[    7135] = 32'h4f738e2a;
    ram_cell[    7136] = 32'h17a39ba2;
    ram_cell[    7137] = 32'h2e44d27c;
    ram_cell[    7138] = 32'he6e753c9;
    ram_cell[    7139] = 32'h1b8aba04;
    ram_cell[    7140] = 32'h0dc9deab;
    ram_cell[    7141] = 32'hb0946a27;
    ram_cell[    7142] = 32'hfcae5912;
    ram_cell[    7143] = 32'hf6092888;
    ram_cell[    7144] = 32'hec328f5b;
    ram_cell[    7145] = 32'he7a5f7c1;
    ram_cell[    7146] = 32'h6bd8acc3;
    ram_cell[    7147] = 32'h89efaa8c;
    ram_cell[    7148] = 32'h51831ce2;
    ram_cell[    7149] = 32'hfc1a377c;
    ram_cell[    7150] = 32'h0c01302e;
    ram_cell[    7151] = 32'h7a77c6d1;
    ram_cell[    7152] = 32'h56ee3f7f;
    ram_cell[    7153] = 32'h3f2e8a7d;
    ram_cell[    7154] = 32'h7eb4d6f6;
    ram_cell[    7155] = 32'hc320e6a2;
    ram_cell[    7156] = 32'hd7c61a32;
    ram_cell[    7157] = 32'h189db376;
    ram_cell[    7158] = 32'h14d8993e;
    ram_cell[    7159] = 32'h69ef6f0c;
    ram_cell[    7160] = 32'h0c280114;
    ram_cell[    7161] = 32'hc4a49a08;
    ram_cell[    7162] = 32'h045e4c38;
    ram_cell[    7163] = 32'h2b9c453a;
    ram_cell[    7164] = 32'h96890186;
    ram_cell[    7165] = 32'h4e3d422a;
    ram_cell[    7166] = 32'h8ced0706;
    ram_cell[    7167] = 32'hf112534b;
    ram_cell[    7168] = 32'h6c84e09b;
    ram_cell[    7169] = 32'had1b13fa;
    ram_cell[    7170] = 32'h56ae6ec2;
    ram_cell[    7171] = 32'h115bd8b2;
    ram_cell[    7172] = 32'he019fa77;
    ram_cell[    7173] = 32'hba662136;
    ram_cell[    7174] = 32'haa5b1c3c;
    ram_cell[    7175] = 32'h3428ea84;
    ram_cell[    7176] = 32'h484cabae;
    ram_cell[    7177] = 32'h8a667749;
    ram_cell[    7178] = 32'hbaad372c;
    ram_cell[    7179] = 32'h31a4d59a;
    ram_cell[    7180] = 32'h5a27fa3e;
    ram_cell[    7181] = 32'h4551d733;
    ram_cell[    7182] = 32'h6b8066e4;
    ram_cell[    7183] = 32'hc0c19543;
    ram_cell[    7184] = 32'hd5506d15;
    ram_cell[    7185] = 32'h633d32e1;
    ram_cell[    7186] = 32'hd65b5789;
    ram_cell[    7187] = 32'h67bfc588;
    ram_cell[    7188] = 32'h96b8ff5b;
    ram_cell[    7189] = 32'h593fa283;
    ram_cell[    7190] = 32'h821f52dd;
    ram_cell[    7191] = 32'ha996e109;
    ram_cell[    7192] = 32'h5439e63b;
    ram_cell[    7193] = 32'hf0d712cd;
    ram_cell[    7194] = 32'heab42387;
    ram_cell[    7195] = 32'h27351475;
    ram_cell[    7196] = 32'h1d37ee45;
    ram_cell[    7197] = 32'h5ace5f38;
    ram_cell[    7198] = 32'he892e0dc;
    ram_cell[    7199] = 32'h3684e8d2;
    ram_cell[    7200] = 32'h28208586;
    ram_cell[    7201] = 32'he7e3fee0;
    ram_cell[    7202] = 32'h0993ddb7;
    ram_cell[    7203] = 32'hcdaf4420;
    ram_cell[    7204] = 32'h375ecd2d;
    ram_cell[    7205] = 32'h3285b6d6;
    ram_cell[    7206] = 32'h0b770cf9;
    ram_cell[    7207] = 32'h305d537f;
    ram_cell[    7208] = 32'h6effdaae;
    ram_cell[    7209] = 32'hc2574752;
    ram_cell[    7210] = 32'h1dc9f962;
    ram_cell[    7211] = 32'hde0af378;
    ram_cell[    7212] = 32'h311ff8de;
    ram_cell[    7213] = 32'h9314db40;
    ram_cell[    7214] = 32'ha2e13a1f;
    ram_cell[    7215] = 32'hdce00ea7;
    ram_cell[    7216] = 32'h2d7d7b23;
    ram_cell[    7217] = 32'ha17104d3;
    ram_cell[    7218] = 32'he36e7a83;
    ram_cell[    7219] = 32'hcc663b59;
    ram_cell[    7220] = 32'h4c92c55c;
    ram_cell[    7221] = 32'hf7224278;
    ram_cell[    7222] = 32'ha0046f5b;
    ram_cell[    7223] = 32'hc4a8aa2c;
    ram_cell[    7224] = 32'hc4900190;
    ram_cell[    7225] = 32'h2fe401ac;
    ram_cell[    7226] = 32'h900787e8;
    ram_cell[    7227] = 32'h5abbbe26;
    ram_cell[    7228] = 32'hcaf05b84;
    ram_cell[    7229] = 32'h3618dd6d;
    ram_cell[    7230] = 32'h315efde7;
    ram_cell[    7231] = 32'h00173d70;
    ram_cell[    7232] = 32'h85997b50;
    ram_cell[    7233] = 32'h60abc938;
    ram_cell[    7234] = 32'hb72e5c4f;
    ram_cell[    7235] = 32'h87c10f24;
    ram_cell[    7236] = 32'h8ba3e05f;
    ram_cell[    7237] = 32'h56bba0e3;
    ram_cell[    7238] = 32'he9c7e785;
    ram_cell[    7239] = 32'h9656e385;
    ram_cell[    7240] = 32'h522d87d9;
    ram_cell[    7241] = 32'ha1a81697;
    ram_cell[    7242] = 32'h7c6e32e9;
    ram_cell[    7243] = 32'h915e7341;
    ram_cell[    7244] = 32'hfdd37c71;
    ram_cell[    7245] = 32'h060c9694;
    ram_cell[    7246] = 32'h12adb3c7;
    ram_cell[    7247] = 32'ha7d51a37;
    ram_cell[    7248] = 32'h85256bbd;
    ram_cell[    7249] = 32'hc1eb9ac1;
    ram_cell[    7250] = 32'h94e7a801;
    ram_cell[    7251] = 32'ha9687a1a;
    ram_cell[    7252] = 32'h62461d55;
    ram_cell[    7253] = 32'h952f17ba;
    ram_cell[    7254] = 32'he6992437;
    ram_cell[    7255] = 32'h4e7adcce;
    ram_cell[    7256] = 32'hff2309ae;
    ram_cell[    7257] = 32'h112ba5da;
    ram_cell[    7258] = 32'hc671a610;
    ram_cell[    7259] = 32'h2124e7aa;
    ram_cell[    7260] = 32'he754d084;
    ram_cell[    7261] = 32'h363a4987;
    ram_cell[    7262] = 32'hd25b0f44;
    ram_cell[    7263] = 32'h7c190e11;
    ram_cell[    7264] = 32'h9ed44085;
    ram_cell[    7265] = 32'hf5174f70;
    ram_cell[    7266] = 32'h2392ca72;
    ram_cell[    7267] = 32'he49f298f;
    ram_cell[    7268] = 32'hb179876f;
    ram_cell[    7269] = 32'h2822c318;
    ram_cell[    7270] = 32'h3d0b24cc;
    ram_cell[    7271] = 32'h579743ba;
    ram_cell[    7272] = 32'h19dde3fe;
    ram_cell[    7273] = 32'h27fa831b;
    ram_cell[    7274] = 32'hdbf2bb05;
    ram_cell[    7275] = 32'h9788c025;
    ram_cell[    7276] = 32'h52b12fe9;
    ram_cell[    7277] = 32'h9b18e56c;
    ram_cell[    7278] = 32'h45765fcb;
    ram_cell[    7279] = 32'h12a3c292;
    ram_cell[    7280] = 32'h1b74e07b;
    ram_cell[    7281] = 32'h218409be;
    ram_cell[    7282] = 32'h2407713a;
    ram_cell[    7283] = 32'hc5b37200;
    ram_cell[    7284] = 32'h1afd1029;
    ram_cell[    7285] = 32'h18ae822e;
    ram_cell[    7286] = 32'h7f45c1c6;
    ram_cell[    7287] = 32'h78d586f4;
    ram_cell[    7288] = 32'h3dc4a75c;
    ram_cell[    7289] = 32'hb2d1c79c;
    ram_cell[    7290] = 32'hedcd4008;
    ram_cell[    7291] = 32'hb641eb5f;
    ram_cell[    7292] = 32'h39ae0bfa;
    ram_cell[    7293] = 32'h1cc7f228;
    ram_cell[    7294] = 32'h4bb9687e;
    ram_cell[    7295] = 32'h3950574f;
    ram_cell[    7296] = 32'hd50c86b5;
    ram_cell[    7297] = 32'ha4f9a157;
    ram_cell[    7298] = 32'h0575db6f;
    ram_cell[    7299] = 32'h830d2d32;
    ram_cell[    7300] = 32'hdf89de0f;
    ram_cell[    7301] = 32'h5cea9542;
    ram_cell[    7302] = 32'h174150d2;
    ram_cell[    7303] = 32'h2e967d74;
    ram_cell[    7304] = 32'h1c3981a2;
    ram_cell[    7305] = 32'hd7bded90;
    ram_cell[    7306] = 32'h596675f2;
    ram_cell[    7307] = 32'hb2e4b81f;
    ram_cell[    7308] = 32'h266c3359;
    ram_cell[    7309] = 32'h07e00df0;
    ram_cell[    7310] = 32'h7f85637d;
    ram_cell[    7311] = 32'h671f4d7d;
    ram_cell[    7312] = 32'hf03fbbb0;
    ram_cell[    7313] = 32'hca3ca870;
    ram_cell[    7314] = 32'h58aaf708;
    ram_cell[    7315] = 32'h4afcef6e;
    ram_cell[    7316] = 32'h39bb9b86;
    ram_cell[    7317] = 32'h10811916;
    ram_cell[    7318] = 32'h5e68df7c;
    ram_cell[    7319] = 32'h8eba8e62;
    ram_cell[    7320] = 32'h9dbc782a;
    ram_cell[    7321] = 32'h2485f252;
    ram_cell[    7322] = 32'h63bacc9c;
    ram_cell[    7323] = 32'h84414c50;
    ram_cell[    7324] = 32'h7aa18f5d;
    ram_cell[    7325] = 32'ha742e593;
    ram_cell[    7326] = 32'h7ae80f64;
    ram_cell[    7327] = 32'hc6a94ba8;
    ram_cell[    7328] = 32'h9b7a851e;
    ram_cell[    7329] = 32'h70cba14d;
    ram_cell[    7330] = 32'h4a36f9bf;
    ram_cell[    7331] = 32'h9e8fe286;
    ram_cell[    7332] = 32'h01524e80;
    ram_cell[    7333] = 32'hc29aa61b;
    ram_cell[    7334] = 32'h4b4bb220;
    ram_cell[    7335] = 32'h3e58962b;
    ram_cell[    7336] = 32'h0c331841;
    ram_cell[    7337] = 32'he5902cef;
    ram_cell[    7338] = 32'h7f29a2d3;
    ram_cell[    7339] = 32'h7dbe8ff4;
    ram_cell[    7340] = 32'hfceaa5f9;
    ram_cell[    7341] = 32'h07c7a58d;
    ram_cell[    7342] = 32'hfd6907ba;
    ram_cell[    7343] = 32'h6b311024;
    ram_cell[    7344] = 32'hecdc2c8b;
    ram_cell[    7345] = 32'hee00649d;
    ram_cell[    7346] = 32'hbf94a24f;
    ram_cell[    7347] = 32'h664305f8;
    ram_cell[    7348] = 32'h59c03134;
    ram_cell[    7349] = 32'hca38310f;
    ram_cell[    7350] = 32'hc8d8c2af;
    ram_cell[    7351] = 32'habf1cd70;
    ram_cell[    7352] = 32'h7902a1b3;
    ram_cell[    7353] = 32'h332f5685;
    ram_cell[    7354] = 32'h1fa2fffb;
    ram_cell[    7355] = 32'hd6b44959;
    ram_cell[    7356] = 32'h095c9ef5;
    ram_cell[    7357] = 32'hda1d6be6;
    ram_cell[    7358] = 32'hb67b1405;
    ram_cell[    7359] = 32'hb7da1c26;
    ram_cell[    7360] = 32'hff4826fb;
    ram_cell[    7361] = 32'h8904df42;
    ram_cell[    7362] = 32'h0264a2c2;
    ram_cell[    7363] = 32'h0e9fda7f;
    ram_cell[    7364] = 32'hb671112a;
    ram_cell[    7365] = 32'h76c47ac4;
    ram_cell[    7366] = 32'h38c38baa;
    ram_cell[    7367] = 32'hd9fcc78b;
    ram_cell[    7368] = 32'h2a46b1f5;
    ram_cell[    7369] = 32'h49600316;
    ram_cell[    7370] = 32'h81d7222b;
    ram_cell[    7371] = 32'hdac5e27b;
    ram_cell[    7372] = 32'h2927b430;
    ram_cell[    7373] = 32'hde4fd839;
    ram_cell[    7374] = 32'h3a84f68d;
    ram_cell[    7375] = 32'hef6debb4;
    ram_cell[    7376] = 32'ha8845b00;
    ram_cell[    7377] = 32'h17741a2a;
    ram_cell[    7378] = 32'ha52446cf;
    ram_cell[    7379] = 32'h0a248e91;
    ram_cell[    7380] = 32'hc44524b5;
    ram_cell[    7381] = 32'he7694ac6;
    ram_cell[    7382] = 32'h96c66a76;
    ram_cell[    7383] = 32'hdd6fea82;
    ram_cell[    7384] = 32'haf2db19a;
    ram_cell[    7385] = 32'h0e64e7ad;
    ram_cell[    7386] = 32'hf0999ed5;
    ram_cell[    7387] = 32'hb9074a71;
    ram_cell[    7388] = 32'hc9b112d2;
    ram_cell[    7389] = 32'he0d8e623;
    ram_cell[    7390] = 32'ha602fb0b;
    ram_cell[    7391] = 32'h53640ba3;
    ram_cell[    7392] = 32'hf57a1235;
    ram_cell[    7393] = 32'h9a61be8b;
    ram_cell[    7394] = 32'h21f166b9;
    ram_cell[    7395] = 32'h450ff70e;
    ram_cell[    7396] = 32'h8e4f60ca;
    ram_cell[    7397] = 32'h6636cd0f;
    ram_cell[    7398] = 32'haa6bb256;
    ram_cell[    7399] = 32'he9766094;
    ram_cell[    7400] = 32'h97278ceb;
    ram_cell[    7401] = 32'h98efaf48;
    ram_cell[    7402] = 32'hba6e8c7c;
    ram_cell[    7403] = 32'hf7c79ac1;
    ram_cell[    7404] = 32'hb5ccbb72;
    ram_cell[    7405] = 32'ha5b6171f;
    ram_cell[    7406] = 32'h1f32d637;
    ram_cell[    7407] = 32'hbf1afb14;
    ram_cell[    7408] = 32'h449c411e;
    ram_cell[    7409] = 32'hbab19c19;
    ram_cell[    7410] = 32'h12ab0acf;
    ram_cell[    7411] = 32'hbc21852f;
    ram_cell[    7412] = 32'h02e29fea;
    ram_cell[    7413] = 32'h27892c49;
    ram_cell[    7414] = 32'h8355f234;
    ram_cell[    7415] = 32'hcddc77da;
    ram_cell[    7416] = 32'hd69307a0;
    ram_cell[    7417] = 32'h181f8853;
    ram_cell[    7418] = 32'haadf3f09;
    ram_cell[    7419] = 32'h8907b007;
    ram_cell[    7420] = 32'hb633ef51;
    ram_cell[    7421] = 32'h12e63e08;
    ram_cell[    7422] = 32'h7369b2fd;
    ram_cell[    7423] = 32'h9b46be39;
    ram_cell[    7424] = 32'h4a2aa89d;
    ram_cell[    7425] = 32'h809f4a96;
    ram_cell[    7426] = 32'h8af0b878;
    ram_cell[    7427] = 32'hd893c9f5;
    ram_cell[    7428] = 32'hb9b23a18;
    ram_cell[    7429] = 32'h335ed7d2;
    ram_cell[    7430] = 32'h4935631b;
    ram_cell[    7431] = 32'h1b09722f;
    ram_cell[    7432] = 32'hd11c3872;
    ram_cell[    7433] = 32'ha224b857;
    ram_cell[    7434] = 32'hcc4e4427;
    ram_cell[    7435] = 32'hb126820c;
    ram_cell[    7436] = 32'hc9732547;
    ram_cell[    7437] = 32'hc4be3b57;
    ram_cell[    7438] = 32'hfc49e811;
    ram_cell[    7439] = 32'hf23764fd;
    ram_cell[    7440] = 32'h43873508;
    ram_cell[    7441] = 32'h355aa1de;
    ram_cell[    7442] = 32'ha469ec67;
    ram_cell[    7443] = 32'h6c5edfe2;
    ram_cell[    7444] = 32'h23965093;
    ram_cell[    7445] = 32'hbfa4a5c1;
    ram_cell[    7446] = 32'hdfc01389;
    ram_cell[    7447] = 32'h9082d2f2;
    ram_cell[    7448] = 32'h1d5c1b04;
    ram_cell[    7449] = 32'h6d65ed90;
    ram_cell[    7450] = 32'h1b44e6f4;
    ram_cell[    7451] = 32'hae719e4e;
    ram_cell[    7452] = 32'h55eae6bf;
    ram_cell[    7453] = 32'h88ea2a35;
    ram_cell[    7454] = 32'hdb377fa2;
    ram_cell[    7455] = 32'ha8fea835;
    ram_cell[    7456] = 32'hdfddcc54;
    ram_cell[    7457] = 32'h8bbc84d0;
    ram_cell[    7458] = 32'hfec16d17;
    ram_cell[    7459] = 32'hcb346ed8;
    ram_cell[    7460] = 32'h0014e89f;
    ram_cell[    7461] = 32'h14e3d68e;
    ram_cell[    7462] = 32'hec28e519;
    ram_cell[    7463] = 32'hc66145b7;
    ram_cell[    7464] = 32'hd0416244;
    ram_cell[    7465] = 32'h1327769e;
    ram_cell[    7466] = 32'h6523e343;
    ram_cell[    7467] = 32'hc1ac17fb;
    ram_cell[    7468] = 32'h98a314d2;
    ram_cell[    7469] = 32'hc2fc2881;
    ram_cell[    7470] = 32'h2e123ce7;
    ram_cell[    7471] = 32'hed7f0f39;
    ram_cell[    7472] = 32'ha0a08f1b;
    ram_cell[    7473] = 32'hc0b4b8ad;
    ram_cell[    7474] = 32'he44504a7;
    ram_cell[    7475] = 32'h9cc97e2c;
    ram_cell[    7476] = 32'ha221f446;
    ram_cell[    7477] = 32'h6d5fa13f;
    ram_cell[    7478] = 32'hc1a22308;
    ram_cell[    7479] = 32'hf389fe7c;
    ram_cell[    7480] = 32'h0b243bbc;
    ram_cell[    7481] = 32'hb66a3d00;
    ram_cell[    7482] = 32'h2f252b16;
    ram_cell[    7483] = 32'hb7147ef1;
    ram_cell[    7484] = 32'hbc8e1948;
    ram_cell[    7485] = 32'h3c69d526;
    ram_cell[    7486] = 32'h29fc2e85;
    ram_cell[    7487] = 32'h33222d10;
    ram_cell[    7488] = 32'h038c9a49;
    ram_cell[    7489] = 32'h3f4a1ff7;
    ram_cell[    7490] = 32'h3f5182a6;
    ram_cell[    7491] = 32'hdd442967;
    ram_cell[    7492] = 32'h207da824;
    ram_cell[    7493] = 32'h95e5357a;
    ram_cell[    7494] = 32'h208f8f48;
    ram_cell[    7495] = 32'h5a947d1e;
    ram_cell[    7496] = 32'hf001b9ab;
    ram_cell[    7497] = 32'h640eef57;
    ram_cell[    7498] = 32'hcfb4224d;
    ram_cell[    7499] = 32'h0d7a10e5;
    ram_cell[    7500] = 32'h6792faa1;
    ram_cell[    7501] = 32'h0259c80a;
    ram_cell[    7502] = 32'hf6638b58;
    ram_cell[    7503] = 32'h6435c0ee;
    ram_cell[    7504] = 32'h7b139c63;
    ram_cell[    7505] = 32'he23164d3;
    ram_cell[    7506] = 32'h97745125;
    ram_cell[    7507] = 32'h279b38fb;
    ram_cell[    7508] = 32'hc7d6ed64;
    ram_cell[    7509] = 32'hcb0fdb54;
    ram_cell[    7510] = 32'h7637bf7a;
    ram_cell[    7511] = 32'h31df8dba;
    ram_cell[    7512] = 32'hb9db4726;
    ram_cell[    7513] = 32'h0b8725f3;
    ram_cell[    7514] = 32'h4253dc06;
    ram_cell[    7515] = 32'h7ee43514;
    ram_cell[    7516] = 32'h4ac8067c;
    ram_cell[    7517] = 32'haeaa317a;
    ram_cell[    7518] = 32'h1ce2ef29;
    ram_cell[    7519] = 32'h09c64b59;
    ram_cell[    7520] = 32'h8eee99dd;
    ram_cell[    7521] = 32'h0a210db2;
    ram_cell[    7522] = 32'he46f0f9e;
    ram_cell[    7523] = 32'h5a91428e;
    ram_cell[    7524] = 32'hdb679e72;
    ram_cell[    7525] = 32'h41e76813;
    ram_cell[    7526] = 32'ha9eaff4b;
    ram_cell[    7527] = 32'h463daa6b;
    ram_cell[    7528] = 32'hf62ed6c5;
    ram_cell[    7529] = 32'h042c93ec;
    ram_cell[    7530] = 32'h7c420766;
    ram_cell[    7531] = 32'hd2c2aaa5;
    ram_cell[    7532] = 32'h984db92d;
    ram_cell[    7533] = 32'hb9975e6d;
    ram_cell[    7534] = 32'he2730bc9;
    ram_cell[    7535] = 32'h0276a01e;
    ram_cell[    7536] = 32'hf1bc0cdd;
    ram_cell[    7537] = 32'h1df73e8e;
    ram_cell[    7538] = 32'h4ccccb60;
    ram_cell[    7539] = 32'h768b0a17;
    ram_cell[    7540] = 32'hcb2d2df8;
    ram_cell[    7541] = 32'h54140820;
    ram_cell[    7542] = 32'h81f53cbe;
    ram_cell[    7543] = 32'h36984ff4;
    ram_cell[    7544] = 32'h9f10c948;
    ram_cell[    7545] = 32'h6a002dd6;
    ram_cell[    7546] = 32'h941ed91c;
    ram_cell[    7547] = 32'hfcc28411;
    ram_cell[    7548] = 32'h13a43300;
    ram_cell[    7549] = 32'he0b435f1;
    ram_cell[    7550] = 32'h6cfe5723;
    ram_cell[    7551] = 32'hc8668adc;
    ram_cell[    7552] = 32'h12a14068;
    ram_cell[    7553] = 32'h10ba9d8a;
    ram_cell[    7554] = 32'hefd894f8;
    ram_cell[    7555] = 32'h3b901b27;
    ram_cell[    7556] = 32'hcae6a128;
    ram_cell[    7557] = 32'h4141b4b5;
    ram_cell[    7558] = 32'he3d3a722;
    ram_cell[    7559] = 32'he3987834;
    ram_cell[    7560] = 32'h5e18fb7d;
    ram_cell[    7561] = 32'ha8e8a82b;
    ram_cell[    7562] = 32'h89c2acdf;
    ram_cell[    7563] = 32'hcaf7300d;
    ram_cell[    7564] = 32'h9df8e08e;
    ram_cell[    7565] = 32'h619092f8;
    ram_cell[    7566] = 32'h90371441;
    ram_cell[    7567] = 32'h460ee907;
    ram_cell[    7568] = 32'h72c8661b;
    ram_cell[    7569] = 32'hfbe274d0;
    ram_cell[    7570] = 32'h3dc9f41a;
    ram_cell[    7571] = 32'h92396a0a;
    ram_cell[    7572] = 32'hff61b25d;
    ram_cell[    7573] = 32'ha7c5f309;
    ram_cell[    7574] = 32'hbdd1518e;
    ram_cell[    7575] = 32'hf00df100;
    ram_cell[    7576] = 32'haaec7e23;
    ram_cell[    7577] = 32'h893256ab;
    ram_cell[    7578] = 32'hfec01994;
    ram_cell[    7579] = 32'h468e886d;
    ram_cell[    7580] = 32'h43af4bec;
    ram_cell[    7581] = 32'hcb9d58c5;
    ram_cell[    7582] = 32'h521a050f;
    ram_cell[    7583] = 32'h0f4a63d1;
    ram_cell[    7584] = 32'h4b9531d6;
    ram_cell[    7585] = 32'h5ee6fff7;
    ram_cell[    7586] = 32'h57097981;
    ram_cell[    7587] = 32'hc8e9efb0;
    ram_cell[    7588] = 32'h80b859e3;
    ram_cell[    7589] = 32'he63b0e1f;
    ram_cell[    7590] = 32'h5d75cde8;
    ram_cell[    7591] = 32'h2e702097;
    ram_cell[    7592] = 32'h0e2f000f;
    ram_cell[    7593] = 32'h32b5918d;
    ram_cell[    7594] = 32'h5eb13de6;
    ram_cell[    7595] = 32'h2088c745;
    ram_cell[    7596] = 32'h9f23d3d8;
    ram_cell[    7597] = 32'h65c8e5c7;
    ram_cell[    7598] = 32'h7e334f6f;
    ram_cell[    7599] = 32'haffa74e7;
    ram_cell[    7600] = 32'h1df307dd;
    ram_cell[    7601] = 32'hefca6c2f;
    ram_cell[    7602] = 32'hfffdbbbb;
    ram_cell[    7603] = 32'h468c9e78;
    ram_cell[    7604] = 32'hbe3a9578;
    ram_cell[    7605] = 32'hf13014c1;
    ram_cell[    7606] = 32'ha9d980f5;
    ram_cell[    7607] = 32'h720ef4e9;
    ram_cell[    7608] = 32'h4c6a7d36;
    ram_cell[    7609] = 32'h2f283376;
    ram_cell[    7610] = 32'h7dfca204;
    ram_cell[    7611] = 32'hb69f9124;
    ram_cell[    7612] = 32'ha597870e;
    ram_cell[    7613] = 32'hc4990418;
    ram_cell[    7614] = 32'hbced8468;
    ram_cell[    7615] = 32'hea55058d;
    ram_cell[    7616] = 32'h24e1955d;
    ram_cell[    7617] = 32'h585c0f22;
    ram_cell[    7618] = 32'h7e55d24a;
    ram_cell[    7619] = 32'h37c65975;
    ram_cell[    7620] = 32'hf0260f2e;
    ram_cell[    7621] = 32'hd8c3393d;
    ram_cell[    7622] = 32'hed74457a;
    ram_cell[    7623] = 32'h4967edc8;
    ram_cell[    7624] = 32'ha694b87f;
    ram_cell[    7625] = 32'hb786cc3f;
    ram_cell[    7626] = 32'h8a796421;
    ram_cell[    7627] = 32'hcb135173;
    ram_cell[    7628] = 32'ha6a0b3cf;
    ram_cell[    7629] = 32'hf7ec2e2e;
    ram_cell[    7630] = 32'hdfbaddee;
    ram_cell[    7631] = 32'h7c0ca11c;
    ram_cell[    7632] = 32'ha6ff9e50;
    ram_cell[    7633] = 32'h52b5d859;
    ram_cell[    7634] = 32'haff0038d;
    ram_cell[    7635] = 32'h6ce9ab1a;
    ram_cell[    7636] = 32'hccff0d36;
    ram_cell[    7637] = 32'hc50e7530;
    ram_cell[    7638] = 32'he9faddcc;
    ram_cell[    7639] = 32'h4515d9fd;
    ram_cell[    7640] = 32'h576ef38e;
    ram_cell[    7641] = 32'h369501d4;
    ram_cell[    7642] = 32'h2542e1b6;
    ram_cell[    7643] = 32'h4da9d84d;
    ram_cell[    7644] = 32'hf097b60e;
    ram_cell[    7645] = 32'h182811b6;
    ram_cell[    7646] = 32'hb0659b88;
    ram_cell[    7647] = 32'h7906b427;
    ram_cell[    7648] = 32'h0739861e;
    ram_cell[    7649] = 32'h3925cb54;
    ram_cell[    7650] = 32'h922dd1cc;
    ram_cell[    7651] = 32'hd35422bc;
    ram_cell[    7652] = 32'h651380a8;
    ram_cell[    7653] = 32'h05e84072;
    ram_cell[    7654] = 32'h3150d946;
    ram_cell[    7655] = 32'hef5c0b12;
    ram_cell[    7656] = 32'hd806e232;
    ram_cell[    7657] = 32'hcc06d101;
    ram_cell[    7658] = 32'h42245279;
    ram_cell[    7659] = 32'h6ba43c77;
    ram_cell[    7660] = 32'hb6d7557a;
    ram_cell[    7661] = 32'hc3ff725d;
    ram_cell[    7662] = 32'h26170bc3;
    ram_cell[    7663] = 32'h3363296c;
    ram_cell[    7664] = 32'hdc7498ef;
    ram_cell[    7665] = 32'h090931da;
    ram_cell[    7666] = 32'h56eb7813;
    ram_cell[    7667] = 32'hbb16f6b7;
    ram_cell[    7668] = 32'h639d1ad0;
    ram_cell[    7669] = 32'hbf932a32;
    ram_cell[    7670] = 32'h7b5b3f38;
    ram_cell[    7671] = 32'h7c8b7220;
    ram_cell[    7672] = 32'h3d0a62c3;
    ram_cell[    7673] = 32'h7a64d7d2;
    ram_cell[    7674] = 32'h3a103bdf;
    ram_cell[    7675] = 32'hbfc1cb0b;
    ram_cell[    7676] = 32'h95cefeac;
    ram_cell[    7677] = 32'h94c8d223;
    ram_cell[    7678] = 32'h212a3bef;
    ram_cell[    7679] = 32'he2f55808;
    ram_cell[    7680] = 32'h593ae988;
    ram_cell[    7681] = 32'hcb4d9e54;
    ram_cell[    7682] = 32'h9c4979ce;
    ram_cell[    7683] = 32'h973c3b3f;
    ram_cell[    7684] = 32'h52f48701;
    ram_cell[    7685] = 32'hfdee7628;
    ram_cell[    7686] = 32'h9c999367;
    ram_cell[    7687] = 32'haab6deb7;
    ram_cell[    7688] = 32'h3fe22b91;
    ram_cell[    7689] = 32'hba3e405a;
    ram_cell[    7690] = 32'h304978cc;
    ram_cell[    7691] = 32'h4d87eb57;
    ram_cell[    7692] = 32'h823fe686;
    ram_cell[    7693] = 32'hd83e4d44;
    ram_cell[    7694] = 32'h2f6ec70c;
    ram_cell[    7695] = 32'hebd26fbf;
    ram_cell[    7696] = 32'h2f10685d;
    ram_cell[    7697] = 32'h2e8733ac;
    ram_cell[    7698] = 32'h327d0d99;
    ram_cell[    7699] = 32'h74643a81;
    ram_cell[    7700] = 32'hae0d7682;
    ram_cell[    7701] = 32'hd67c77ba;
    ram_cell[    7702] = 32'hb12f131e;
    ram_cell[    7703] = 32'h0d90f14a;
    ram_cell[    7704] = 32'h5d0b9b92;
    ram_cell[    7705] = 32'h7af930e3;
    ram_cell[    7706] = 32'h4447219d;
    ram_cell[    7707] = 32'h729f9c1e;
    ram_cell[    7708] = 32'he9c35adc;
    ram_cell[    7709] = 32'h291e5eb4;
    ram_cell[    7710] = 32'hd1ab0045;
    ram_cell[    7711] = 32'he42c37fe;
    ram_cell[    7712] = 32'h79d0e591;
    ram_cell[    7713] = 32'h60a5d949;
    ram_cell[    7714] = 32'h9a5f0c34;
    ram_cell[    7715] = 32'hfd6ae6a0;
    ram_cell[    7716] = 32'h2ebb6b25;
    ram_cell[    7717] = 32'hb756ffb8;
    ram_cell[    7718] = 32'h325a1c30;
    ram_cell[    7719] = 32'hea57cbbc;
    ram_cell[    7720] = 32'hca4bec8d;
    ram_cell[    7721] = 32'habdca063;
    ram_cell[    7722] = 32'h10882f65;
    ram_cell[    7723] = 32'h8a9d5f28;
    ram_cell[    7724] = 32'h070d1c3d;
    ram_cell[    7725] = 32'he0b4852c;
    ram_cell[    7726] = 32'hdba77c53;
    ram_cell[    7727] = 32'h9ded4580;
    ram_cell[    7728] = 32'hfd8e3a80;
    ram_cell[    7729] = 32'hccc19489;
    ram_cell[    7730] = 32'h73c3e10e;
    ram_cell[    7731] = 32'h817852e2;
    ram_cell[    7732] = 32'hc46aea03;
    ram_cell[    7733] = 32'hf5e2bb62;
    ram_cell[    7734] = 32'hbbabf5b9;
    ram_cell[    7735] = 32'h31038110;
    ram_cell[    7736] = 32'hec19322b;
    ram_cell[    7737] = 32'h3a7facf8;
    ram_cell[    7738] = 32'hfc58da7b;
    ram_cell[    7739] = 32'h570237bc;
    ram_cell[    7740] = 32'hba572d94;
    ram_cell[    7741] = 32'h0604a9d8;
    ram_cell[    7742] = 32'h9a5064f1;
    ram_cell[    7743] = 32'hb1af5fc6;
    ram_cell[    7744] = 32'h4b86b5e6;
    ram_cell[    7745] = 32'h288e4e10;
    ram_cell[    7746] = 32'h1d80cb4e;
    ram_cell[    7747] = 32'h1049dcac;
    ram_cell[    7748] = 32'h729fc19a;
    ram_cell[    7749] = 32'he48ebd53;
    ram_cell[    7750] = 32'h19e46451;
    ram_cell[    7751] = 32'hd22b408f;
    ram_cell[    7752] = 32'he767ce0a;
    ram_cell[    7753] = 32'h49c1c9f8;
    ram_cell[    7754] = 32'h1a127e79;
    ram_cell[    7755] = 32'h1ade79b2;
    ram_cell[    7756] = 32'hdc099c09;
    ram_cell[    7757] = 32'h2f73fdc3;
    ram_cell[    7758] = 32'hb29a5424;
    ram_cell[    7759] = 32'h4e7d6960;
    ram_cell[    7760] = 32'hca6eed58;
    ram_cell[    7761] = 32'he0d09325;
    ram_cell[    7762] = 32'h633102b7;
    ram_cell[    7763] = 32'h838db057;
    ram_cell[    7764] = 32'hea28bd0d;
    ram_cell[    7765] = 32'hb4fd2ced;
    ram_cell[    7766] = 32'h3c095b34;
    ram_cell[    7767] = 32'hc56c250b;
    ram_cell[    7768] = 32'h18ff63bd;
    ram_cell[    7769] = 32'he51533ae;
    ram_cell[    7770] = 32'h3410574c;
    ram_cell[    7771] = 32'h73922403;
    ram_cell[    7772] = 32'hbbaec82a;
    ram_cell[    7773] = 32'haed91a80;
    ram_cell[    7774] = 32'h6954d8d1;
    ram_cell[    7775] = 32'h9583e079;
    ram_cell[    7776] = 32'h7f029ed9;
    ram_cell[    7777] = 32'h43dfc4f0;
    ram_cell[    7778] = 32'h4c686ccc;
    ram_cell[    7779] = 32'h0dffc46b;
    ram_cell[    7780] = 32'h9d48e875;
    ram_cell[    7781] = 32'hcf19c385;
    ram_cell[    7782] = 32'hce6af28f;
    ram_cell[    7783] = 32'hc7fdd589;
    ram_cell[    7784] = 32'h63e32384;
    ram_cell[    7785] = 32'hda5ac9a6;
    ram_cell[    7786] = 32'h16f25278;
    ram_cell[    7787] = 32'h505f172e;
    ram_cell[    7788] = 32'h96265a30;
    ram_cell[    7789] = 32'hdb6153dc;
    ram_cell[    7790] = 32'h5bfdb65d;
    ram_cell[    7791] = 32'hab0c2643;
    ram_cell[    7792] = 32'h22752574;
    ram_cell[    7793] = 32'ha04378f5;
    ram_cell[    7794] = 32'hb9d8f564;
    ram_cell[    7795] = 32'hcc81c0e8;
    ram_cell[    7796] = 32'h7b49b7cf;
    ram_cell[    7797] = 32'h2a97987c;
    ram_cell[    7798] = 32'h00c3f26b;
    ram_cell[    7799] = 32'he5cc6579;
    ram_cell[    7800] = 32'h803ca3dd;
    ram_cell[    7801] = 32'h20d7b060;
    ram_cell[    7802] = 32'hb58470c7;
    ram_cell[    7803] = 32'hcdbd5ea5;
    ram_cell[    7804] = 32'h40296326;
    ram_cell[    7805] = 32'he1c3e26b;
    ram_cell[    7806] = 32'h4c1ef5d8;
    ram_cell[    7807] = 32'hc99e011a;
    ram_cell[    7808] = 32'hc8c48593;
    ram_cell[    7809] = 32'h92ed6b81;
    ram_cell[    7810] = 32'hb67da5e5;
    ram_cell[    7811] = 32'h4d82fa1c;
    ram_cell[    7812] = 32'he1365cae;
    ram_cell[    7813] = 32'hd9819bb9;
    ram_cell[    7814] = 32'h10c46744;
    ram_cell[    7815] = 32'heeda0102;
    ram_cell[    7816] = 32'h9be694fa;
    ram_cell[    7817] = 32'h9ab4e1e6;
    ram_cell[    7818] = 32'h12bb7b9b;
    ram_cell[    7819] = 32'hf09da6c6;
    ram_cell[    7820] = 32'h39e681ba;
    ram_cell[    7821] = 32'h00bc00de;
    ram_cell[    7822] = 32'h5dea5bdd;
    ram_cell[    7823] = 32'hd6ce5306;
    ram_cell[    7824] = 32'hc0ccae7b;
    ram_cell[    7825] = 32'hc034c09a;
    ram_cell[    7826] = 32'h2f58e837;
    ram_cell[    7827] = 32'h09e1d951;
    ram_cell[    7828] = 32'h2f1c0e6d;
    ram_cell[    7829] = 32'hfcd03260;
    ram_cell[    7830] = 32'h1758b21b;
    ram_cell[    7831] = 32'h535eedc2;
    ram_cell[    7832] = 32'h07651b51;
    ram_cell[    7833] = 32'hd99df975;
    ram_cell[    7834] = 32'h51e58020;
    ram_cell[    7835] = 32'ha780a4a5;
    ram_cell[    7836] = 32'hfbd21747;
    ram_cell[    7837] = 32'h8afaabf9;
    ram_cell[    7838] = 32'hf7f20250;
    ram_cell[    7839] = 32'hc2133a48;
    ram_cell[    7840] = 32'hd91adee5;
    ram_cell[    7841] = 32'h0cdc8178;
    ram_cell[    7842] = 32'h1d0ce439;
    ram_cell[    7843] = 32'ha9150810;
    ram_cell[    7844] = 32'h76c3c048;
    ram_cell[    7845] = 32'hcb326dfe;
    ram_cell[    7846] = 32'h06e8d816;
    ram_cell[    7847] = 32'h83bfd401;
    ram_cell[    7848] = 32'h86b65a36;
    ram_cell[    7849] = 32'h9c67aabf;
    ram_cell[    7850] = 32'h4174d877;
    ram_cell[    7851] = 32'h87fc8673;
    ram_cell[    7852] = 32'h9ca5a206;
    ram_cell[    7853] = 32'h35f39aba;
    ram_cell[    7854] = 32'h361df859;
    ram_cell[    7855] = 32'h030b988a;
    ram_cell[    7856] = 32'hfd8580cf;
    ram_cell[    7857] = 32'h5fa02324;
    ram_cell[    7858] = 32'h3b16bc5d;
    ram_cell[    7859] = 32'h2db8cd87;
    ram_cell[    7860] = 32'hb1f93314;
    ram_cell[    7861] = 32'h3edacab6;
    ram_cell[    7862] = 32'h9b9e638e;
    ram_cell[    7863] = 32'hb22d5c70;
    ram_cell[    7864] = 32'h0e83caa8;
    ram_cell[    7865] = 32'had947803;
    ram_cell[    7866] = 32'hdeddad97;
    ram_cell[    7867] = 32'h4fcbfe96;
    ram_cell[    7868] = 32'hb9366f6b;
    ram_cell[    7869] = 32'h68b3e1e5;
    ram_cell[    7870] = 32'h68203e86;
    ram_cell[    7871] = 32'hb08c379c;
    ram_cell[    7872] = 32'h38dd51bc;
    ram_cell[    7873] = 32'h815fa132;
    ram_cell[    7874] = 32'h690c85d1;
    ram_cell[    7875] = 32'he6ed263e;
    ram_cell[    7876] = 32'h540363bd;
    ram_cell[    7877] = 32'h6b841c7e;
    ram_cell[    7878] = 32'h4685c3a8;
    ram_cell[    7879] = 32'hb2d4a072;
    ram_cell[    7880] = 32'hf1f4664d;
    ram_cell[    7881] = 32'h484e14bd;
    ram_cell[    7882] = 32'h51b2fb26;
    ram_cell[    7883] = 32'hb77234b9;
    ram_cell[    7884] = 32'h63537506;
    ram_cell[    7885] = 32'h9e0d61e5;
    ram_cell[    7886] = 32'hfa4085ad;
    ram_cell[    7887] = 32'h2b42be9f;
    ram_cell[    7888] = 32'hf12c2954;
    ram_cell[    7889] = 32'h55c78c17;
    ram_cell[    7890] = 32'h33f5315e;
    ram_cell[    7891] = 32'hce9ca4a7;
    ram_cell[    7892] = 32'h1b59f7a5;
    ram_cell[    7893] = 32'h020f27e9;
    ram_cell[    7894] = 32'hacbc44ea;
    ram_cell[    7895] = 32'h727a956c;
    ram_cell[    7896] = 32'h756419d7;
    ram_cell[    7897] = 32'h1421d80a;
    ram_cell[    7898] = 32'he6e63ce8;
    ram_cell[    7899] = 32'h90cb167c;
    ram_cell[    7900] = 32'h43f97b6c;
    ram_cell[    7901] = 32'ha98656f1;
    ram_cell[    7902] = 32'h16d626bb;
    ram_cell[    7903] = 32'h4f3f78b9;
    ram_cell[    7904] = 32'h231899a7;
    ram_cell[    7905] = 32'h5d7936ef;
    ram_cell[    7906] = 32'h233bbfe1;
    ram_cell[    7907] = 32'h68b51737;
    ram_cell[    7908] = 32'hfa3be5a7;
    ram_cell[    7909] = 32'haa29f89f;
    ram_cell[    7910] = 32'h86913fd5;
    ram_cell[    7911] = 32'hf29d63d4;
    ram_cell[    7912] = 32'hc79db493;
    ram_cell[    7913] = 32'h3cd40055;
    ram_cell[    7914] = 32'h5d60134e;
    ram_cell[    7915] = 32'h08307abe;
    ram_cell[    7916] = 32'h4fd810b2;
    ram_cell[    7917] = 32'hefa93bc5;
    ram_cell[    7918] = 32'h5fc8d5e2;
    ram_cell[    7919] = 32'h62a24362;
    ram_cell[    7920] = 32'hdccd2726;
    ram_cell[    7921] = 32'h00defdaa;
    ram_cell[    7922] = 32'h95a83f87;
    ram_cell[    7923] = 32'ha2523012;
    ram_cell[    7924] = 32'h5f57e132;
    ram_cell[    7925] = 32'hcd657528;
    ram_cell[    7926] = 32'h8a87f19c;
    ram_cell[    7927] = 32'h76c0c120;
    ram_cell[    7928] = 32'h8944eeec;
    ram_cell[    7929] = 32'h1e5e8e14;
    ram_cell[    7930] = 32'h5889bd3c;
    ram_cell[    7931] = 32'h28f0ef84;
    ram_cell[    7932] = 32'hf02eef11;
    ram_cell[    7933] = 32'h4ae73304;
    ram_cell[    7934] = 32'h395d4b38;
    ram_cell[    7935] = 32'hb15d5afb;
    ram_cell[    7936] = 32'h48f07290;
    ram_cell[    7937] = 32'h4ce07300;
    ram_cell[    7938] = 32'ha479bd87;
    ram_cell[    7939] = 32'hf0dfa3a5;
    ram_cell[    7940] = 32'hb264d046;
    ram_cell[    7941] = 32'heb38240d;
    ram_cell[    7942] = 32'ha018f362;
    ram_cell[    7943] = 32'h89a4a047;
    ram_cell[    7944] = 32'h160c8179;
    ram_cell[    7945] = 32'h551a35a0;
    ram_cell[    7946] = 32'h5e5ece6d;
    ram_cell[    7947] = 32'h1c11d522;
    ram_cell[    7948] = 32'ha69c8dbc;
    ram_cell[    7949] = 32'h77649443;
    ram_cell[    7950] = 32'hc1d48149;
    ram_cell[    7951] = 32'h27bfcecd;
    ram_cell[    7952] = 32'h5bc5a128;
    ram_cell[    7953] = 32'h7180b42a;
    ram_cell[    7954] = 32'h842a7333;
    ram_cell[    7955] = 32'h8066ed67;
    ram_cell[    7956] = 32'hb626d14f;
    ram_cell[    7957] = 32'h507f96cc;
    ram_cell[    7958] = 32'h6a3b35eb;
    ram_cell[    7959] = 32'h8bc96696;
    ram_cell[    7960] = 32'hba3ab3dc;
    ram_cell[    7961] = 32'h7c7faf46;
    ram_cell[    7962] = 32'h51a81fbf;
    ram_cell[    7963] = 32'hfd46aadc;
    ram_cell[    7964] = 32'hc6a82d84;
    ram_cell[    7965] = 32'hdf484da7;
    ram_cell[    7966] = 32'h48cb66a3;
    ram_cell[    7967] = 32'h7fbae357;
    ram_cell[    7968] = 32'h44a3c74a;
    ram_cell[    7969] = 32'he98c980c;
    ram_cell[    7970] = 32'hc9782597;
    ram_cell[    7971] = 32'ha4577787;
    ram_cell[    7972] = 32'hc9984e34;
    ram_cell[    7973] = 32'h9c74091f;
    ram_cell[    7974] = 32'h2c882a40;
    ram_cell[    7975] = 32'hb57bac09;
    ram_cell[    7976] = 32'h332c2e0e;
    ram_cell[    7977] = 32'h28da90ba;
    ram_cell[    7978] = 32'h46fb3c76;
    ram_cell[    7979] = 32'h25572997;
    ram_cell[    7980] = 32'h7ca05855;
    ram_cell[    7981] = 32'ha5806394;
    ram_cell[    7982] = 32'hb355bfeb;
    ram_cell[    7983] = 32'he5c1ee4c;
    ram_cell[    7984] = 32'h3e5ae292;
    ram_cell[    7985] = 32'h96440bcc;
    ram_cell[    7986] = 32'hbe89cdc5;
    ram_cell[    7987] = 32'h14611a4a;
    ram_cell[    7988] = 32'hd22d1528;
    ram_cell[    7989] = 32'hc884e6e9;
    ram_cell[    7990] = 32'hfe8e190b;
    ram_cell[    7991] = 32'h9dab60fa;
    ram_cell[    7992] = 32'hac7453e3;
    ram_cell[    7993] = 32'hee3c6235;
    ram_cell[    7994] = 32'hd579ddbe;
    ram_cell[    7995] = 32'hbdd4e775;
    ram_cell[    7996] = 32'h5eca73b5;
    ram_cell[    7997] = 32'h57ee79b1;
    ram_cell[    7998] = 32'h8c18a890;
    ram_cell[    7999] = 32'h66d9ecbc;
    ram_cell[    8000] = 32'hcd1bffae;
    ram_cell[    8001] = 32'h1369c9f6;
    ram_cell[    8002] = 32'h12026e94;
    ram_cell[    8003] = 32'h35aa7701;
    ram_cell[    8004] = 32'h0bf0a095;
    ram_cell[    8005] = 32'h5b18209b;
    ram_cell[    8006] = 32'h003d6dd7;
    ram_cell[    8007] = 32'hd9d67644;
    ram_cell[    8008] = 32'hc1e9fc6e;
    ram_cell[    8009] = 32'h4da07180;
    ram_cell[    8010] = 32'h321c7d4c;
    ram_cell[    8011] = 32'h18ba9bf9;
    ram_cell[    8012] = 32'hf2e23805;
    ram_cell[    8013] = 32'h1cb69aef;
    ram_cell[    8014] = 32'h0a242d3f;
    ram_cell[    8015] = 32'h0f1b8921;
    ram_cell[    8016] = 32'h057cac10;
    ram_cell[    8017] = 32'hc6b8ad7b;
    ram_cell[    8018] = 32'h284c9f49;
    ram_cell[    8019] = 32'h2f19ecc9;
    ram_cell[    8020] = 32'h9b2b1bf9;
    ram_cell[    8021] = 32'h7bcd508b;
    ram_cell[    8022] = 32'hf28659f3;
    ram_cell[    8023] = 32'h21d832bc;
    ram_cell[    8024] = 32'hfbae51dd;
    ram_cell[    8025] = 32'h44dbd0db;
    ram_cell[    8026] = 32'hf338dee9;
    ram_cell[    8027] = 32'h47149a2f;
    ram_cell[    8028] = 32'h95bdd93b;
    ram_cell[    8029] = 32'hcece4831;
    ram_cell[    8030] = 32'h598879b2;
    ram_cell[    8031] = 32'h0199bf8c;
    ram_cell[    8032] = 32'h22c55d79;
    ram_cell[    8033] = 32'hcbf53396;
    ram_cell[    8034] = 32'hf2ccd67f;
    ram_cell[    8035] = 32'h298dcc49;
    ram_cell[    8036] = 32'h91a30978;
    ram_cell[    8037] = 32'hc254cd12;
    ram_cell[    8038] = 32'h4fd76eff;
    ram_cell[    8039] = 32'h412bb6b6;
    ram_cell[    8040] = 32'haba18570;
    ram_cell[    8041] = 32'h1f0f7a3b;
    ram_cell[    8042] = 32'h59c8699c;
    ram_cell[    8043] = 32'h8433dc32;
    ram_cell[    8044] = 32'h747a1143;
    ram_cell[    8045] = 32'h9f7ad27b;
    ram_cell[    8046] = 32'ha0009be8;
    ram_cell[    8047] = 32'h02fa14b7;
    ram_cell[    8048] = 32'h4ee6622b;
    ram_cell[    8049] = 32'haef80a8b;
    ram_cell[    8050] = 32'he0313ae1;
    ram_cell[    8051] = 32'h3f5ae570;
    ram_cell[    8052] = 32'h8db6bcba;
    ram_cell[    8053] = 32'hca8e1a87;
    ram_cell[    8054] = 32'h4a52b970;
    ram_cell[    8055] = 32'h0509f6bf;
    ram_cell[    8056] = 32'hb913c30f;
    ram_cell[    8057] = 32'h824d7db8;
    ram_cell[    8058] = 32'h5ee7f94e;
    ram_cell[    8059] = 32'hd07820cd;
    ram_cell[    8060] = 32'h28ca1307;
    ram_cell[    8061] = 32'h6d1b9565;
    ram_cell[    8062] = 32'h5fc4d00b;
    ram_cell[    8063] = 32'h77da9195;
    ram_cell[    8064] = 32'h90993462;
    ram_cell[    8065] = 32'hfae6f2dc;
    ram_cell[    8066] = 32'h73d3537a;
    ram_cell[    8067] = 32'h0c4889a0;
    ram_cell[    8068] = 32'h43661af4;
    ram_cell[    8069] = 32'h37700e8b;
    ram_cell[    8070] = 32'hb8b26547;
    ram_cell[    8071] = 32'hcf8f0202;
    ram_cell[    8072] = 32'he580aab6;
    ram_cell[    8073] = 32'ha9177719;
    ram_cell[    8074] = 32'h7cd05965;
    ram_cell[    8075] = 32'hb8de5d48;
    ram_cell[    8076] = 32'haaee18a0;
    ram_cell[    8077] = 32'hfc166b79;
    ram_cell[    8078] = 32'h816e7c5f;
    ram_cell[    8079] = 32'hd175ff70;
    ram_cell[    8080] = 32'h3ec8f76e;
    ram_cell[    8081] = 32'h83cf56e2;
    ram_cell[    8082] = 32'h490cabcb;
    ram_cell[    8083] = 32'h638b9119;
    ram_cell[    8084] = 32'h6c3b7f20;
    ram_cell[    8085] = 32'hb5683630;
    ram_cell[    8086] = 32'hec88b799;
    ram_cell[    8087] = 32'h0b8de5c2;
    ram_cell[    8088] = 32'h49860c69;
    ram_cell[    8089] = 32'h536472f5;
    ram_cell[    8090] = 32'h375a6422;
    ram_cell[    8091] = 32'h3bb828ef;
    ram_cell[    8092] = 32'hb71a283e;
    ram_cell[    8093] = 32'hb6231e6f;
    ram_cell[    8094] = 32'haa2d2382;
    ram_cell[    8095] = 32'habe4485f;
    ram_cell[    8096] = 32'hb3e8dba5;
    ram_cell[    8097] = 32'h5665624a;
    ram_cell[    8098] = 32'hb933094b;
    ram_cell[    8099] = 32'h2215cca5;
    ram_cell[    8100] = 32'hf377d1fe;
    ram_cell[    8101] = 32'h4bdbf5b8;
    ram_cell[    8102] = 32'hd631e0ee;
    ram_cell[    8103] = 32'h6a0ae99a;
    ram_cell[    8104] = 32'hd6313bc4;
    ram_cell[    8105] = 32'h9fa86354;
    ram_cell[    8106] = 32'h4c6eeeb9;
    ram_cell[    8107] = 32'h04188ec3;
    ram_cell[    8108] = 32'h69d42ed5;
    ram_cell[    8109] = 32'h09603834;
    ram_cell[    8110] = 32'h59c6de7b;
    ram_cell[    8111] = 32'h21c99c9e;
    ram_cell[    8112] = 32'h16ad6856;
    ram_cell[    8113] = 32'h5f2d95e3;
    ram_cell[    8114] = 32'hcb03474a;
    ram_cell[    8115] = 32'hf1b4be83;
    ram_cell[    8116] = 32'h3e7b84e3;
    ram_cell[    8117] = 32'h7e8a0b7b;
    ram_cell[    8118] = 32'had9ddfa3;
    ram_cell[    8119] = 32'hf52d426d;
    ram_cell[    8120] = 32'hbd7ea0aa;
    ram_cell[    8121] = 32'h93f940bb;
    ram_cell[    8122] = 32'hd22d762d;
    ram_cell[    8123] = 32'h2508a610;
    ram_cell[    8124] = 32'h24715b39;
    ram_cell[    8125] = 32'hae7b40e2;
    ram_cell[    8126] = 32'h7c9fe79c;
    ram_cell[    8127] = 32'h8cf2c910;
    ram_cell[    8128] = 32'hf98d095f;
    ram_cell[    8129] = 32'hd377ff3d;
    ram_cell[    8130] = 32'h4091779b;
    ram_cell[    8131] = 32'hed0b3377;
    ram_cell[    8132] = 32'h0320acec;
    ram_cell[    8133] = 32'h945a1bef;
    ram_cell[    8134] = 32'hbe2df55e;
    ram_cell[    8135] = 32'hb4f0ac6c;
    ram_cell[    8136] = 32'h92e97550;
    ram_cell[    8137] = 32'h4564142e;
    ram_cell[    8138] = 32'h3c0cc861;
    ram_cell[    8139] = 32'hf75d437e;
    ram_cell[    8140] = 32'h6fe26f62;
    ram_cell[    8141] = 32'hb389151f;
    ram_cell[    8142] = 32'hb4b77d67;
    ram_cell[    8143] = 32'hf5685e4b;
    ram_cell[    8144] = 32'h1f771550;
    ram_cell[    8145] = 32'hc3707115;
    ram_cell[    8146] = 32'ha7ed369d;
    ram_cell[    8147] = 32'h57efd84b;
    ram_cell[    8148] = 32'hccf7f4aa;
    ram_cell[    8149] = 32'h50fcd888;
    ram_cell[    8150] = 32'heb1bd5a0;
    ram_cell[    8151] = 32'hc45a0a91;
    ram_cell[    8152] = 32'hf35ace71;
    ram_cell[    8153] = 32'h37636c95;
    ram_cell[    8154] = 32'hcd73ab45;
    ram_cell[    8155] = 32'h6bbb40ed;
    ram_cell[    8156] = 32'ha9441bf5;
    ram_cell[    8157] = 32'h11fb4325;
    ram_cell[    8158] = 32'h9997327f;
    ram_cell[    8159] = 32'hd4616036;
    ram_cell[    8160] = 32'h1540d058;
    ram_cell[    8161] = 32'h1f4ef342;
    ram_cell[    8162] = 32'hb169a5a5;
    ram_cell[    8163] = 32'h27c9c044;
    ram_cell[    8164] = 32'h5a0e471e;
    ram_cell[    8165] = 32'he94de44e;
    ram_cell[    8166] = 32'ha726012b;
    ram_cell[    8167] = 32'hcf6d08f4;
    ram_cell[    8168] = 32'he878ed3b;
    ram_cell[    8169] = 32'h16dab8da;
    ram_cell[    8170] = 32'h4812093e;
    ram_cell[    8171] = 32'h03199597;
    ram_cell[    8172] = 32'he2cb76aa;
    ram_cell[    8173] = 32'hbb01d72f;
    ram_cell[    8174] = 32'h71a7c7fa;
    ram_cell[    8175] = 32'hb8fca666;
    ram_cell[    8176] = 32'ha2cb4f0d;
    ram_cell[    8177] = 32'h4e2bd0e7;
    ram_cell[    8178] = 32'h825adae2;
    ram_cell[    8179] = 32'h60c8216f;
    ram_cell[    8180] = 32'hdf17b783;
    ram_cell[    8181] = 32'h4d82bb5c;
    ram_cell[    8182] = 32'h33f265aa;
    ram_cell[    8183] = 32'hd42ae31f;
    ram_cell[    8184] = 32'hd0cf8e85;
    ram_cell[    8185] = 32'hfa082dc6;
    ram_cell[    8186] = 32'hbf9369d5;
    ram_cell[    8187] = 32'h6853a41d;
    ram_cell[    8188] = 32'h54415c53;
    ram_cell[    8189] = 32'h93a053ca;
    ram_cell[    8190] = 32'he0aba610;
    ram_cell[    8191] = 32'h236e034a;
    // src matrix B
    ram_cell[    8192] = 32'h411c8100;
    ram_cell[    8193] = 32'h5b3d97a5;
    ram_cell[    8194] = 32'hdd9dd40b;
    ram_cell[    8195] = 32'h0e3bca67;
    ram_cell[    8196] = 32'h981a6adf;
    ram_cell[    8197] = 32'hafb3ae16;
    ram_cell[    8198] = 32'h5e5fec53;
    ram_cell[    8199] = 32'h2afe5905;
    ram_cell[    8200] = 32'h275a164c;
    ram_cell[    8201] = 32'had649d06;
    ram_cell[    8202] = 32'h8b0d6a6a;
    ram_cell[    8203] = 32'h883bad6c;
    ram_cell[    8204] = 32'h967f4336;
    ram_cell[    8205] = 32'hcd4a8ba3;
    ram_cell[    8206] = 32'h9e8dc0a5;
    ram_cell[    8207] = 32'hce6ff457;
    ram_cell[    8208] = 32'h4813cec0;
    ram_cell[    8209] = 32'h8a24b10a;
    ram_cell[    8210] = 32'h854eb781;
    ram_cell[    8211] = 32'hce1d4086;
    ram_cell[    8212] = 32'he650a215;
    ram_cell[    8213] = 32'hfbfd8b79;
    ram_cell[    8214] = 32'h4a8ca789;
    ram_cell[    8215] = 32'he36e713b;
    ram_cell[    8216] = 32'h99fa4173;
    ram_cell[    8217] = 32'h481e3af6;
    ram_cell[    8218] = 32'h6bd78c2a;
    ram_cell[    8219] = 32'h6927fdcf;
    ram_cell[    8220] = 32'h19ad58c7;
    ram_cell[    8221] = 32'h2dab6789;
    ram_cell[    8222] = 32'hf5079046;
    ram_cell[    8223] = 32'h2e258aa6;
    ram_cell[    8224] = 32'h7cda57dc;
    ram_cell[    8225] = 32'ha1e0eb27;
    ram_cell[    8226] = 32'h3860dbde;
    ram_cell[    8227] = 32'hbb90535b;
    ram_cell[    8228] = 32'h07dff07c;
    ram_cell[    8229] = 32'hdff5dbdd;
    ram_cell[    8230] = 32'hec9eafc2;
    ram_cell[    8231] = 32'h0bd97491;
    ram_cell[    8232] = 32'h12dbe793;
    ram_cell[    8233] = 32'h11f15b20;
    ram_cell[    8234] = 32'h0a901899;
    ram_cell[    8235] = 32'h98aac8fa;
    ram_cell[    8236] = 32'hf0de71b5;
    ram_cell[    8237] = 32'hd3409cd0;
    ram_cell[    8238] = 32'h8fba2ce8;
    ram_cell[    8239] = 32'hbaf9d5ca;
    ram_cell[    8240] = 32'he6673f96;
    ram_cell[    8241] = 32'he59133d3;
    ram_cell[    8242] = 32'hc6ffc816;
    ram_cell[    8243] = 32'hbb515693;
    ram_cell[    8244] = 32'h8b952008;
    ram_cell[    8245] = 32'h96c8189b;
    ram_cell[    8246] = 32'hf965c47d;
    ram_cell[    8247] = 32'h4b42c50d;
    ram_cell[    8248] = 32'h4cdfcf35;
    ram_cell[    8249] = 32'h3eabab50;
    ram_cell[    8250] = 32'heda678b8;
    ram_cell[    8251] = 32'h52d83006;
    ram_cell[    8252] = 32'h9d25ae11;
    ram_cell[    8253] = 32'h64c85c48;
    ram_cell[    8254] = 32'h651774e5;
    ram_cell[    8255] = 32'h1c62061d;
    ram_cell[    8256] = 32'hc2aab0cf;
    ram_cell[    8257] = 32'hac2c82cd;
    ram_cell[    8258] = 32'he9c9cbf3;
    ram_cell[    8259] = 32'h88d93c37;
    ram_cell[    8260] = 32'h0ff41cd5;
    ram_cell[    8261] = 32'hea15f414;
    ram_cell[    8262] = 32'h9d355b7e;
    ram_cell[    8263] = 32'h6626bdc1;
    ram_cell[    8264] = 32'h8fcfc86a;
    ram_cell[    8265] = 32'hbeeed9b8;
    ram_cell[    8266] = 32'hc6b95937;
    ram_cell[    8267] = 32'h5ce4059e;
    ram_cell[    8268] = 32'hb73bd69c;
    ram_cell[    8269] = 32'h777aa43e;
    ram_cell[    8270] = 32'h13603a08;
    ram_cell[    8271] = 32'h1ed9238c;
    ram_cell[    8272] = 32'h5acc7f5b;
    ram_cell[    8273] = 32'h26364f11;
    ram_cell[    8274] = 32'h0916200e;
    ram_cell[    8275] = 32'hc3cf67fa;
    ram_cell[    8276] = 32'hc89178f9;
    ram_cell[    8277] = 32'h36bc6519;
    ram_cell[    8278] = 32'h9314e72b;
    ram_cell[    8279] = 32'h86f178e6;
    ram_cell[    8280] = 32'h16f40763;
    ram_cell[    8281] = 32'h08049775;
    ram_cell[    8282] = 32'h3896ac98;
    ram_cell[    8283] = 32'hb4908ae5;
    ram_cell[    8284] = 32'h8e50f16a;
    ram_cell[    8285] = 32'hc3606cea;
    ram_cell[    8286] = 32'ha0f06017;
    ram_cell[    8287] = 32'h898b0a54;
    ram_cell[    8288] = 32'h9171be8a;
    ram_cell[    8289] = 32'h4a32c6b7;
    ram_cell[    8290] = 32'h0aa6f2c6;
    ram_cell[    8291] = 32'h306f2422;
    ram_cell[    8292] = 32'he96e96a7;
    ram_cell[    8293] = 32'hfdfb658d;
    ram_cell[    8294] = 32'hc8b2df33;
    ram_cell[    8295] = 32'h23006834;
    ram_cell[    8296] = 32'h8a9caa60;
    ram_cell[    8297] = 32'hc9056a8e;
    ram_cell[    8298] = 32'h687c6244;
    ram_cell[    8299] = 32'h7e23e0c6;
    ram_cell[    8300] = 32'h3c09cf88;
    ram_cell[    8301] = 32'hea77dec9;
    ram_cell[    8302] = 32'hacac7ab9;
    ram_cell[    8303] = 32'hba39e87c;
    ram_cell[    8304] = 32'heb67c997;
    ram_cell[    8305] = 32'h4f38f8bc;
    ram_cell[    8306] = 32'h09afd5f8;
    ram_cell[    8307] = 32'h68b4a9be;
    ram_cell[    8308] = 32'hba62ad12;
    ram_cell[    8309] = 32'hbd0589d3;
    ram_cell[    8310] = 32'h6231b366;
    ram_cell[    8311] = 32'hbdda5be6;
    ram_cell[    8312] = 32'hf381af1a;
    ram_cell[    8313] = 32'hb0e81b68;
    ram_cell[    8314] = 32'h14c686ac;
    ram_cell[    8315] = 32'h55be7139;
    ram_cell[    8316] = 32'h981092bd;
    ram_cell[    8317] = 32'h92c5574d;
    ram_cell[    8318] = 32'hc314b8b6;
    ram_cell[    8319] = 32'hf487a8bf;
    ram_cell[    8320] = 32'h6a024764;
    ram_cell[    8321] = 32'h8d1799f7;
    ram_cell[    8322] = 32'h713229be;
    ram_cell[    8323] = 32'h9781dca2;
    ram_cell[    8324] = 32'hd9b9eaad;
    ram_cell[    8325] = 32'h6f22b624;
    ram_cell[    8326] = 32'hb3f3306e;
    ram_cell[    8327] = 32'hd126fd81;
    ram_cell[    8328] = 32'hc8e7cc0a;
    ram_cell[    8329] = 32'hbb3a1784;
    ram_cell[    8330] = 32'hee921ec7;
    ram_cell[    8331] = 32'hc7ba0efa;
    ram_cell[    8332] = 32'h0b61526a;
    ram_cell[    8333] = 32'h5dc746b0;
    ram_cell[    8334] = 32'hf1e81a2b;
    ram_cell[    8335] = 32'h065048f5;
    ram_cell[    8336] = 32'h48000a26;
    ram_cell[    8337] = 32'h1a6e199c;
    ram_cell[    8338] = 32'hfe4f54e8;
    ram_cell[    8339] = 32'h2937e7a9;
    ram_cell[    8340] = 32'hb118e932;
    ram_cell[    8341] = 32'hbba7de45;
    ram_cell[    8342] = 32'h50993572;
    ram_cell[    8343] = 32'h93749f39;
    ram_cell[    8344] = 32'h151dfb6e;
    ram_cell[    8345] = 32'hc5bcfee0;
    ram_cell[    8346] = 32'he9be73c5;
    ram_cell[    8347] = 32'h9cf7fa4d;
    ram_cell[    8348] = 32'he5ea3eb3;
    ram_cell[    8349] = 32'h354e73af;
    ram_cell[    8350] = 32'h9839f34f;
    ram_cell[    8351] = 32'h52cc9bb9;
    ram_cell[    8352] = 32'h8d037c95;
    ram_cell[    8353] = 32'hd4d7ce97;
    ram_cell[    8354] = 32'h68bc58f6;
    ram_cell[    8355] = 32'hff22ba22;
    ram_cell[    8356] = 32'h4d8d5d49;
    ram_cell[    8357] = 32'h126a22ba;
    ram_cell[    8358] = 32'hbfcd7c0a;
    ram_cell[    8359] = 32'he20e6911;
    ram_cell[    8360] = 32'h42940c3f;
    ram_cell[    8361] = 32'h5f86e0be;
    ram_cell[    8362] = 32'h5149fb8b;
    ram_cell[    8363] = 32'h3ec41000;
    ram_cell[    8364] = 32'h5259bf73;
    ram_cell[    8365] = 32'h8333a9c1;
    ram_cell[    8366] = 32'hda82a6d9;
    ram_cell[    8367] = 32'hee4ce46e;
    ram_cell[    8368] = 32'h7a761956;
    ram_cell[    8369] = 32'h2ea77587;
    ram_cell[    8370] = 32'he28edd79;
    ram_cell[    8371] = 32'h6e6e9abf;
    ram_cell[    8372] = 32'h0eae8c36;
    ram_cell[    8373] = 32'hbc70614b;
    ram_cell[    8374] = 32'hd471a3a0;
    ram_cell[    8375] = 32'h60daa928;
    ram_cell[    8376] = 32'h0fe70b11;
    ram_cell[    8377] = 32'h0d6a53b6;
    ram_cell[    8378] = 32'hf44747a8;
    ram_cell[    8379] = 32'hf3eb8466;
    ram_cell[    8380] = 32'hf948a43a;
    ram_cell[    8381] = 32'ha1b9ba66;
    ram_cell[    8382] = 32'h9c1473c4;
    ram_cell[    8383] = 32'h45926c17;
    ram_cell[    8384] = 32'h66a2d773;
    ram_cell[    8385] = 32'hc79bf7dc;
    ram_cell[    8386] = 32'hfc8f302f;
    ram_cell[    8387] = 32'ha8ed6124;
    ram_cell[    8388] = 32'hfe466ebd;
    ram_cell[    8389] = 32'h4027bc46;
    ram_cell[    8390] = 32'h39c49a35;
    ram_cell[    8391] = 32'hca36ee5f;
    ram_cell[    8392] = 32'hf0719eeb;
    ram_cell[    8393] = 32'h932dea09;
    ram_cell[    8394] = 32'ha388e55b;
    ram_cell[    8395] = 32'h187a6d92;
    ram_cell[    8396] = 32'h785c641f;
    ram_cell[    8397] = 32'h39c683af;
    ram_cell[    8398] = 32'h25936844;
    ram_cell[    8399] = 32'h08bf6857;
    ram_cell[    8400] = 32'h60bc4ae5;
    ram_cell[    8401] = 32'hfdde38ea;
    ram_cell[    8402] = 32'h84a083dc;
    ram_cell[    8403] = 32'h3bdfd75a;
    ram_cell[    8404] = 32'h98936761;
    ram_cell[    8405] = 32'hf3bccbc2;
    ram_cell[    8406] = 32'h21a8da53;
    ram_cell[    8407] = 32'hdf97e988;
    ram_cell[    8408] = 32'ha32cc773;
    ram_cell[    8409] = 32'hd9912215;
    ram_cell[    8410] = 32'h54c2b26d;
    ram_cell[    8411] = 32'hbf10db78;
    ram_cell[    8412] = 32'h422b8d1e;
    ram_cell[    8413] = 32'ha82e2745;
    ram_cell[    8414] = 32'h022e1957;
    ram_cell[    8415] = 32'hb7a236b3;
    ram_cell[    8416] = 32'h5e02c16c;
    ram_cell[    8417] = 32'hf471eedc;
    ram_cell[    8418] = 32'h7f9b9bb3;
    ram_cell[    8419] = 32'h79f5b74e;
    ram_cell[    8420] = 32'h778ecf2c;
    ram_cell[    8421] = 32'ha431bed8;
    ram_cell[    8422] = 32'ha35522d2;
    ram_cell[    8423] = 32'h01067a1d;
    ram_cell[    8424] = 32'h05602cb9;
    ram_cell[    8425] = 32'h67a644dd;
    ram_cell[    8426] = 32'h56b08545;
    ram_cell[    8427] = 32'hd2fcb1c6;
    ram_cell[    8428] = 32'hbb744fdf;
    ram_cell[    8429] = 32'h94b6a081;
    ram_cell[    8430] = 32'hf9063352;
    ram_cell[    8431] = 32'h6471889f;
    ram_cell[    8432] = 32'hf6b94e21;
    ram_cell[    8433] = 32'hb971ff1d;
    ram_cell[    8434] = 32'h6a5193a0;
    ram_cell[    8435] = 32'hd3f4d343;
    ram_cell[    8436] = 32'hcef4f664;
    ram_cell[    8437] = 32'haf96cff0;
    ram_cell[    8438] = 32'hdf726dde;
    ram_cell[    8439] = 32'h87f2a4f0;
    ram_cell[    8440] = 32'h027a0e0e;
    ram_cell[    8441] = 32'he7d96dfc;
    ram_cell[    8442] = 32'h62bdf62c;
    ram_cell[    8443] = 32'ha316c842;
    ram_cell[    8444] = 32'h8b9b64d0;
    ram_cell[    8445] = 32'hd85b254d;
    ram_cell[    8446] = 32'hbfa0c1d3;
    ram_cell[    8447] = 32'hcf02f6af;
    ram_cell[    8448] = 32'h985f6bd7;
    ram_cell[    8449] = 32'hc92d026c;
    ram_cell[    8450] = 32'h390a9f2b;
    ram_cell[    8451] = 32'hf776185c;
    ram_cell[    8452] = 32'h0ce435e5;
    ram_cell[    8453] = 32'h129ea001;
    ram_cell[    8454] = 32'hc885c38d;
    ram_cell[    8455] = 32'hd6aaa6d2;
    ram_cell[    8456] = 32'h1a86caaf;
    ram_cell[    8457] = 32'h79bbeae5;
    ram_cell[    8458] = 32'hbc9dc9d3;
    ram_cell[    8459] = 32'h933971c8;
    ram_cell[    8460] = 32'h41322dd6;
    ram_cell[    8461] = 32'haacf8030;
    ram_cell[    8462] = 32'h3b5504a9;
    ram_cell[    8463] = 32'hc897b564;
    ram_cell[    8464] = 32'h9c7816c2;
    ram_cell[    8465] = 32'ha30b8b96;
    ram_cell[    8466] = 32'hf99c8076;
    ram_cell[    8467] = 32'h54930fbd;
    ram_cell[    8468] = 32'h22abb59f;
    ram_cell[    8469] = 32'hc24b0a72;
    ram_cell[    8470] = 32'hb33aace1;
    ram_cell[    8471] = 32'hfe3470c9;
    ram_cell[    8472] = 32'h7b9360d0;
    ram_cell[    8473] = 32'h14473964;
    ram_cell[    8474] = 32'h451d90ed;
    ram_cell[    8475] = 32'hbe485c76;
    ram_cell[    8476] = 32'h078091f5;
    ram_cell[    8477] = 32'h4270f8e3;
    ram_cell[    8478] = 32'h30417462;
    ram_cell[    8479] = 32'h618372dc;
    ram_cell[    8480] = 32'hf9d9b1f7;
    ram_cell[    8481] = 32'hb5469a17;
    ram_cell[    8482] = 32'h6141cf6c;
    ram_cell[    8483] = 32'hd89f96cc;
    ram_cell[    8484] = 32'h91dbc144;
    ram_cell[    8485] = 32'h0fe1b995;
    ram_cell[    8486] = 32'h889ef89e;
    ram_cell[    8487] = 32'h5194df51;
    ram_cell[    8488] = 32'h3b6f1343;
    ram_cell[    8489] = 32'hfc2990d6;
    ram_cell[    8490] = 32'ha3955ff7;
    ram_cell[    8491] = 32'hca94ccb8;
    ram_cell[    8492] = 32'h923bd63d;
    ram_cell[    8493] = 32'hcc203ee7;
    ram_cell[    8494] = 32'hd3e7657f;
    ram_cell[    8495] = 32'haf669557;
    ram_cell[    8496] = 32'hc4449039;
    ram_cell[    8497] = 32'h28310c3c;
    ram_cell[    8498] = 32'hd7925ef1;
    ram_cell[    8499] = 32'h88fc0672;
    ram_cell[    8500] = 32'h8319a73e;
    ram_cell[    8501] = 32'h3d5460c9;
    ram_cell[    8502] = 32'hb43992e1;
    ram_cell[    8503] = 32'he7dcf6db;
    ram_cell[    8504] = 32'h0046492f;
    ram_cell[    8505] = 32'h0b12c533;
    ram_cell[    8506] = 32'hac7c0342;
    ram_cell[    8507] = 32'hc0436d5f;
    ram_cell[    8508] = 32'h8437a79b;
    ram_cell[    8509] = 32'h3c75b545;
    ram_cell[    8510] = 32'hdc7e88d1;
    ram_cell[    8511] = 32'hd9470150;
    ram_cell[    8512] = 32'h9b5c5eed;
    ram_cell[    8513] = 32'he8f8415a;
    ram_cell[    8514] = 32'h0a85e964;
    ram_cell[    8515] = 32'h2250b60e;
    ram_cell[    8516] = 32'h8975088b;
    ram_cell[    8517] = 32'hb84bdd2a;
    ram_cell[    8518] = 32'h27ba9867;
    ram_cell[    8519] = 32'h8ce70288;
    ram_cell[    8520] = 32'h0e58b62a;
    ram_cell[    8521] = 32'h2361e781;
    ram_cell[    8522] = 32'heb407f12;
    ram_cell[    8523] = 32'h01904778;
    ram_cell[    8524] = 32'h75e10237;
    ram_cell[    8525] = 32'h77ec5f7d;
    ram_cell[    8526] = 32'h684af65f;
    ram_cell[    8527] = 32'h50b6623e;
    ram_cell[    8528] = 32'hbc7ec7bd;
    ram_cell[    8529] = 32'h0ee6bb5e;
    ram_cell[    8530] = 32'hf3bf340f;
    ram_cell[    8531] = 32'ha9aaf30b;
    ram_cell[    8532] = 32'hfe83b894;
    ram_cell[    8533] = 32'h4ee08cb5;
    ram_cell[    8534] = 32'h77adf927;
    ram_cell[    8535] = 32'h279ec957;
    ram_cell[    8536] = 32'hf1a939fc;
    ram_cell[    8537] = 32'he3d93406;
    ram_cell[    8538] = 32'h21548380;
    ram_cell[    8539] = 32'ha6ba6779;
    ram_cell[    8540] = 32'he601ae3a;
    ram_cell[    8541] = 32'hc0e707d4;
    ram_cell[    8542] = 32'hc9443ba1;
    ram_cell[    8543] = 32'h5392d73e;
    ram_cell[    8544] = 32'hb5e74c99;
    ram_cell[    8545] = 32'ha1575a2b;
    ram_cell[    8546] = 32'he49f22ee;
    ram_cell[    8547] = 32'h18ea5881;
    ram_cell[    8548] = 32'h800ab28e;
    ram_cell[    8549] = 32'hcdcd7f83;
    ram_cell[    8550] = 32'hb08bc115;
    ram_cell[    8551] = 32'h1bb81618;
    ram_cell[    8552] = 32'h9f0f7e88;
    ram_cell[    8553] = 32'h54a6144e;
    ram_cell[    8554] = 32'h0dc6520d;
    ram_cell[    8555] = 32'h2be37bea;
    ram_cell[    8556] = 32'h749d3c64;
    ram_cell[    8557] = 32'h7f2cd58a;
    ram_cell[    8558] = 32'h26294e5b;
    ram_cell[    8559] = 32'h7884b2bb;
    ram_cell[    8560] = 32'ha8c2e2fc;
    ram_cell[    8561] = 32'hcb91c6cb;
    ram_cell[    8562] = 32'h9475f48d;
    ram_cell[    8563] = 32'hca42b881;
    ram_cell[    8564] = 32'h4051b44e;
    ram_cell[    8565] = 32'h1c151ffa;
    ram_cell[    8566] = 32'hedcf26f9;
    ram_cell[    8567] = 32'h3366b42e;
    ram_cell[    8568] = 32'hc2814f7f;
    ram_cell[    8569] = 32'haaa4ced1;
    ram_cell[    8570] = 32'h49ec06c6;
    ram_cell[    8571] = 32'h4d085fca;
    ram_cell[    8572] = 32'hba5807c3;
    ram_cell[    8573] = 32'h16c1c32c;
    ram_cell[    8574] = 32'h5c047423;
    ram_cell[    8575] = 32'h7e34e831;
    ram_cell[    8576] = 32'ha5e519c0;
    ram_cell[    8577] = 32'h57835975;
    ram_cell[    8578] = 32'h4aca87f4;
    ram_cell[    8579] = 32'h7e0e214d;
    ram_cell[    8580] = 32'hddf6a90a;
    ram_cell[    8581] = 32'hdc8eebcb;
    ram_cell[    8582] = 32'hc529c45b;
    ram_cell[    8583] = 32'h305ce2da;
    ram_cell[    8584] = 32'h1c0ba55e;
    ram_cell[    8585] = 32'h77530017;
    ram_cell[    8586] = 32'ha7550086;
    ram_cell[    8587] = 32'h3cc1d6bf;
    ram_cell[    8588] = 32'h6c451e5a;
    ram_cell[    8589] = 32'hd46284f6;
    ram_cell[    8590] = 32'h6d5b5154;
    ram_cell[    8591] = 32'h2a1cdf83;
    ram_cell[    8592] = 32'haf0071fa;
    ram_cell[    8593] = 32'h0f0a73c1;
    ram_cell[    8594] = 32'h79231733;
    ram_cell[    8595] = 32'h370eccfc;
    ram_cell[    8596] = 32'h6e192000;
    ram_cell[    8597] = 32'hdd59a2e7;
    ram_cell[    8598] = 32'h70eace41;
    ram_cell[    8599] = 32'hba8a4985;
    ram_cell[    8600] = 32'h0b703e27;
    ram_cell[    8601] = 32'hd41453ec;
    ram_cell[    8602] = 32'h66f5d722;
    ram_cell[    8603] = 32'h6c5c515a;
    ram_cell[    8604] = 32'h1fbf21f2;
    ram_cell[    8605] = 32'h4885f6b6;
    ram_cell[    8606] = 32'hc831144f;
    ram_cell[    8607] = 32'h8a315596;
    ram_cell[    8608] = 32'hc12537fd;
    ram_cell[    8609] = 32'h3edaa6ec;
    ram_cell[    8610] = 32'hf98aa358;
    ram_cell[    8611] = 32'h86a554fa;
    ram_cell[    8612] = 32'h766604eb;
    ram_cell[    8613] = 32'he2a99291;
    ram_cell[    8614] = 32'hd905f803;
    ram_cell[    8615] = 32'h5fb70f1a;
    ram_cell[    8616] = 32'h12aa81d4;
    ram_cell[    8617] = 32'h2be2dd42;
    ram_cell[    8618] = 32'h88089939;
    ram_cell[    8619] = 32'hb09656ad;
    ram_cell[    8620] = 32'h2b67c760;
    ram_cell[    8621] = 32'h6c14690f;
    ram_cell[    8622] = 32'hf11c7e0c;
    ram_cell[    8623] = 32'h4a9e2d70;
    ram_cell[    8624] = 32'h4f88bed7;
    ram_cell[    8625] = 32'h1b4626c8;
    ram_cell[    8626] = 32'h43cfa726;
    ram_cell[    8627] = 32'h462e1860;
    ram_cell[    8628] = 32'hba82439f;
    ram_cell[    8629] = 32'h08059fa0;
    ram_cell[    8630] = 32'hcb45608c;
    ram_cell[    8631] = 32'h5ba83640;
    ram_cell[    8632] = 32'h5f60af66;
    ram_cell[    8633] = 32'hbef847ac;
    ram_cell[    8634] = 32'h5c391af8;
    ram_cell[    8635] = 32'h3c57621f;
    ram_cell[    8636] = 32'h57df5268;
    ram_cell[    8637] = 32'hfef16325;
    ram_cell[    8638] = 32'h5fc999ee;
    ram_cell[    8639] = 32'hadf98f2d;
    ram_cell[    8640] = 32'h27665f3b;
    ram_cell[    8641] = 32'hd36e314c;
    ram_cell[    8642] = 32'hef99d16c;
    ram_cell[    8643] = 32'h851b5418;
    ram_cell[    8644] = 32'h0b238a53;
    ram_cell[    8645] = 32'hd9822f3e;
    ram_cell[    8646] = 32'h61d5c5d2;
    ram_cell[    8647] = 32'h2a8a60bf;
    ram_cell[    8648] = 32'hbf764dd2;
    ram_cell[    8649] = 32'h1a1dc192;
    ram_cell[    8650] = 32'h1c81b75a;
    ram_cell[    8651] = 32'h75b5a21f;
    ram_cell[    8652] = 32'h271a0753;
    ram_cell[    8653] = 32'hea5f2102;
    ram_cell[    8654] = 32'h0432f663;
    ram_cell[    8655] = 32'hd27e4e00;
    ram_cell[    8656] = 32'h6c020933;
    ram_cell[    8657] = 32'h24e82da3;
    ram_cell[    8658] = 32'h328e93ad;
    ram_cell[    8659] = 32'h0466abd9;
    ram_cell[    8660] = 32'hd33c8788;
    ram_cell[    8661] = 32'h5f6e9bda;
    ram_cell[    8662] = 32'h1e6c8194;
    ram_cell[    8663] = 32'hd2315128;
    ram_cell[    8664] = 32'hd73cc430;
    ram_cell[    8665] = 32'h06310324;
    ram_cell[    8666] = 32'h6d03360d;
    ram_cell[    8667] = 32'h4b831770;
    ram_cell[    8668] = 32'hbd1d1016;
    ram_cell[    8669] = 32'h0e1d01fb;
    ram_cell[    8670] = 32'h4b82c21c;
    ram_cell[    8671] = 32'h18e2dea1;
    ram_cell[    8672] = 32'h060b23c8;
    ram_cell[    8673] = 32'ha7a62559;
    ram_cell[    8674] = 32'h06fe698c;
    ram_cell[    8675] = 32'h91769f8a;
    ram_cell[    8676] = 32'h835d80cc;
    ram_cell[    8677] = 32'h8546053a;
    ram_cell[    8678] = 32'h562fedcf;
    ram_cell[    8679] = 32'h5536b28e;
    ram_cell[    8680] = 32'h84b2532e;
    ram_cell[    8681] = 32'h45eeb27f;
    ram_cell[    8682] = 32'h9eadb4f2;
    ram_cell[    8683] = 32'haf72cb2c;
    ram_cell[    8684] = 32'hed3e7130;
    ram_cell[    8685] = 32'h8ddb3888;
    ram_cell[    8686] = 32'h4f70c1fb;
    ram_cell[    8687] = 32'h8e82bbfd;
    ram_cell[    8688] = 32'h1fc1e038;
    ram_cell[    8689] = 32'hf78f1f13;
    ram_cell[    8690] = 32'h266e4d98;
    ram_cell[    8691] = 32'h1b761fee;
    ram_cell[    8692] = 32'h4e5634b9;
    ram_cell[    8693] = 32'hd8a7e771;
    ram_cell[    8694] = 32'hdd9a5be3;
    ram_cell[    8695] = 32'he17f9594;
    ram_cell[    8696] = 32'h63aeed80;
    ram_cell[    8697] = 32'h5b8027cf;
    ram_cell[    8698] = 32'h881af2af;
    ram_cell[    8699] = 32'hb3f1e8ad;
    ram_cell[    8700] = 32'h7e6ebfb5;
    ram_cell[    8701] = 32'hcd09fcac;
    ram_cell[    8702] = 32'h043f9e47;
    ram_cell[    8703] = 32'h8dcf908c;
    ram_cell[    8704] = 32'h9d5991c2;
    ram_cell[    8705] = 32'h83a35883;
    ram_cell[    8706] = 32'h77e58a57;
    ram_cell[    8707] = 32'h52a4b18b;
    ram_cell[    8708] = 32'hcdfb788d;
    ram_cell[    8709] = 32'h16329cd3;
    ram_cell[    8710] = 32'h75e1195d;
    ram_cell[    8711] = 32'hbd137a14;
    ram_cell[    8712] = 32'hec3eb0e4;
    ram_cell[    8713] = 32'h0bbe16b8;
    ram_cell[    8714] = 32'hd91f2a93;
    ram_cell[    8715] = 32'hb007b730;
    ram_cell[    8716] = 32'h1a81e0ee;
    ram_cell[    8717] = 32'hb461270b;
    ram_cell[    8718] = 32'h8b92be77;
    ram_cell[    8719] = 32'hd25167b7;
    ram_cell[    8720] = 32'hfe24c3fc;
    ram_cell[    8721] = 32'h5b1be014;
    ram_cell[    8722] = 32'h13e7f777;
    ram_cell[    8723] = 32'hd21f676f;
    ram_cell[    8724] = 32'h83d2121f;
    ram_cell[    8725] = 32'h09a977b7;
    ram_cell[    8726] = 32'h779920c0;
    ram_cell[    8727] = 32'h603af766;
    ram_cell[    8728] = 32'hbbda061d;
    ram_cell[    8729] = 32'hd721dfa7;
    ram_cell[    8730] = 32'h1795c252;
    ram_cell[    8731] = 32'ha5ce440d;
    ram_cell[    8732] = 32'hd7175b92;
    ram_cell[    8733] = 32'h1be59b9e;
    ram_cell[    8734] = 32'h0d9380b9;
    ram_cell[    8735] = 32'h41ae7505;
    ram_cell[    8736] = 32'hdc856032;
    ram_cell[    8737] = 32'h2d9ffadf;
    ram_cell[    8738] = 32'h955ec16a;
    ram_cell[    8739] = 32'hd2d49113;
    ram_cell[    8740] = 32'h105195e8;
    ram_cell[    8741] = 32'hdf033045;
    ram_cell[    8742] = 32'he19923e5;
    ram_cell[    8743] = 32'hf8ddee23;
    ram_cell[    8744] = 32'hb8b79d66;
    ram_cell[    8745] = 32'hd5f93ae8;
    ram_cell[    8746] = 32'h52b319ff;
    ram_cell[    8747] = 32'hbc8d668e;
    ram_cell[    8748] = 32'h01d0dd90;
    ram_cell[    8749] = 32'h4b2d26b9;
    ram_cell[    8750] = 32'hbd18b8e9;
    ram_cell[    8751] = 32'hb7ea9f20;
    ram_cell[    8752] = 32'h11e66025;
    ram_cell[    8753] = 32'h933d9454;
    ram_cell[    8754] = 32'hce8fdee6;
    ram_cell[    8755] = 32'h471b039b;
    ram_cell[    8756] = 32'h0f408736;
    ram_cell[    8757] = 32'hf1e31efa;
    ram_cell[    8758] = 32'h64907213;
    ram_cell[    8759] = 32'h0f6e17d1;
    ram_cell[    8760] = 32'hc9ab0431;
    ram_cell[    8761] = 32'h04befb1d;
    ram_cell[    8762] = 32'h645a8c03;
    ram_cell[    8763] = 32'ha40e0144;
    ram_cell[    8764] = 32'h58f2c706;
    ram_cell[    8765] = 32'h0fa83cee;
    ram_cell[    8766] = 32'h1977e46c;
    ram_cell[    8767] = 32'hd8b66ca8;
    ram_cell[    8768] = 32'h1eb91b8b;
    ram_cell[    8769] = 32'hc8012610;
    ram_cell[    8770] = 32'he8ca7981;
    ram_cell[    8771] = 32'h963ab07a;
    ram_cell[    8772] = 32'hce1a6178;
    ram_cell[    8773] = 32'h9a84536e;
    ram_cell[    8774] = 32'h448acc9b;
    ram_cell[    8775] = 32'hc1d06d59;
    ram_cell[    8776] = 32'h83c6e8ad;
    ram_cell[    8777] = 32'hc28caa73;
    ram_cell[    8778] = 32'h5f75fded;
    ram_cell[    8779] = 32'h20fee1d5;
    ram_cell[    8780] = 32'hda7c393e;
    ram_cell[    8781] = 32'h0ffd62cd;
    ram_cell[    8782] = 32'h61f483de;
    ram_cell[    8783] = 32'h1d389567;
    ram_cell[    8784] = 32'h52d94c98;
    ram_cell[    8785] = 32'h20acc043;
    ram_cell[    8786] = 32'hf9b4172e;
    ram_cell[    8787] = 32'h13b3667c;
    ram_cell[    8788] = 32'ha1e65c53;
    ram_cell[    8789] = 32'h2641459f;
    ram_cell[    8790] = 32'he4c5b46b;
    ram_cell[    8791] = 32'h364ec811;
    ram_cell[    8792] = 32'h622a31c2;
    ram_cell[    8793] = 32'heff01931;
    ram_cell[    8794] = 32'he44178f8;
    ram_cell[    8795] = 32'h73091b5f;
    ram_cell[    8796] = 32'he0232f25;
    ram_cell[    8797] = 32'h6a08c7de;
    ram_cell[    8798] = 32'h194f26ab;
    ram_cell[    8799] = 32'h37f5b7f9;
    ram_cell[    8800] = 32'hae918973;
    ram_cell[    8801] = 32'h0eea90c1;
    ram_cell[    8802] = 32'h9a4b0587;
    ram_cell[    8803] = 32'h47485de4;
    ram_cell[    8804] = 32'h4249daaa;
    ram_cell[    8805] = 32'h402527d3;
    ram_cell[    8806] = 32'h676bffe2;
    ram_cell[    8807] = 32'he8964602;
    ram_cell[    8808] = 32'h4f8a2dae;
    ram_cell[    8809] = 32'hbacf5027;
    ram_cell[    8810] = 32'h55f7bb71;
    ram_cell[    8811] = 32'hb9b92b8f;
    ram_cell[    8812] = 32'hbe63163f;
    ram_cell[    8813] = 32'h71bc9735;
    ram_cell[    8814] = 32'hf0b845b6;
    ram_cell[    8815] = 32'hd9d06b58;
    ram_cell[    8816] = 32'h08c643af;
    ram_cell[    8817] = 32'h2996e6e1;
    ram_cell[    8818] = 32'h3d3a232f;
    ram_cell[    8819] = 32'h16146d3d;
    ram_cell[    8820] = 32'h487dc510;
    ram_cell[    8821] = 32'h4893c820;
    ram_cell[    8822] = 32'h017260dd;
    ram_cell[    8823] = 32'hd9835724;
    ram_cell[    8824] = 32'hfbd1e2ac;
    ram_cell[    8825] = 32'he6a5590d;
    ram_cell[    8826] = 32'h1e5631d0;
    ram_cell[    8827] = 32'h52b2e054;
    ram_cell[    8828] = 32'h99a44203;
    ram_cell[    8829] = 32'hc3441fda;
    ram_cell[    8830] = 32'he84aef05;
    ram_cell[    8831] = 32'hf681b799;
    ram_cell[    8832] = 32'h8ed1c105;
    ram_cell[    8833] = 32'h00b2c2c0;
    ram_cell[    8834] = 32'hdc4061bf;
    ram_cell[    8835] = 32'hc8db15e4;
    ram_cell[    8836] = 32'h7c05bc63;
    ram_cell[    8837] = 32'h32d0bafe;
    ram_cell[    8838] = 32'h6b92467d;
    ram_cell[    8839] = 32'h9a4ae787;
    ram_cell[    8840] = 32'hba5e1b24;
    ram_cell[    8841] = 32'hbe33135f;
    ram_cell[    8842] = 32'h529654c9;
    ram_cell[    8843] = 32'he1baf72e;
    ram_cell[    8844] = 32'h43ea3dc1;
    ram_cell[    8845] = 32'h6beb6b80;
    ram_cell[    8846] = 32'h486a291e;
    ram_cell[    8847] = 32'h61a08b15;
    ram_cell[    8848] = 32'hf2467c5d;
    ram_cell[    8849] = 32'hd16c9a8b;
    ram_cell[    8850] = 32'h790cd33e;
    ram_cell[    8851] = 32'h4827c050;
    ram_cell[    8852] = 32'h04f0702e;
    ram_cell[    8853] = 32'hd4fa0ae6;
    ram_cell[    8854] = 32'hbdcf182d;
    ram_cell[    8855] = 32'hef053804;
    ram_cell[    8856] = 32'h1b2e8cbc;
    ram_cell[    8857] = 32'h6c29c688;
    ram_cell[    8858] = 32'hf0a00e2f;
    ram_cell[    8859] = 32'h319788cb;
    ram_cell[    8860] = 32'hb350fbd2;
    ram_cell[    8861] = 32'h073861e0;
    ram_cell[    8862] = 32'h32d02f47;
    ram_cell[    8863] = 32'haa5c7009;
    ram_cell[    8864] = 32'h6b9c6c7b;
    ram_cell[    8865] = 32'h684247b3;
    ram_cell[    8866] = 32'hd660bb48;
    ram_cell[    8867] = 32'h65661341;
    ram_cell[    8868] = 32'h769dcf30;
    ram_cell[    8869] = 32'hd877f7c8;
    ram_cell[    8870] = 32'h8e96b783;
    ram_cell[    8871] = 32'h45c4135e;
    ram_cell[    8872] = 32'h87e8e0a9;
    ram_cell[    8873] = 32'h6fcd152e;
    ram_cell[    8874] = 32'hd35c3968;
    ram_cell[    8875] = 32'h9ff89427;
    ram_cell[    8876] = 32'h65253d76;
    ram_cell[    8877] = 32'h94674f2b;
    ram_cell[    8878] = 32'h2b8a3ccb;
    ram_cell[    8879] = 32'h17ab20ac;
    ram_cell[    8880] = 32'h8d4bc4ec;
    ram_cell[    8881] = 32'h00602db3;
    ram_cell[    8882] = 32'ha0ddddbe;
    ram_cell[    8883] = 32'h58804c11;
    ram_cell[    8884] = 32'h2fbd5550;
    ram_cell[    8885] = 32'hc852ae23;
    ram_cell[    8886] = 32'hc2f7694a;
    ram_cell[    8887] = 32'h5420dc37;
    ram_cell[    8888] = 32'hd77e9d91;
    ram_cell[    8889] = 32'h144a729c;
    ram_cell[    8890] = 32'h9847f25d;
    ram_cell[    8891] = 32'hb68a48de;
    ram_cell[    8892] = 32'h111bad0d;
    ram_cell[    8893] = 32'h685bf9da;
    ram_cell[    8894] = 32'hf65cc74d;
    ram_cell[    8895] = 32'hf29f19fa;
    ram_cell[    8896] = 32'h342f13c2;
    ram_cell[    8897] = 32'h6df57caf;
    ram_cell[    8898] = 32'hfbea6aab;
    ram_cell[    8899] = 32'h5f2843d7;
    ram_cell[    8900] = 32'he709a612;
    ram_cell[    8901] = 32'h1ee447ec;
    ram_cell[    8902] = 32'h0741b397;
    ram_cell[    8903] = 32'h82baadbf;
    ram_cell[    8904] = 32'he41ab71e;
    ram_cell[    8905] = 32'h562fea9b;
    ram_cell[    8906] = 32'h7358187f;
    ram_cell[    8907] = 32'h7273ccff;
    ram_cell[    8908] = 32'h0aeb6bf3;
    ram_cell[    8909] = 32'h684ce6c4;
    ram_cell[    8910] = 32'he8da21da;
    ram_cell[    8911] = 32'hd513a9e9;
    ram_cell[    8912] = 32'h77c69976;
    ram_cell[    8913] = 32'h0d85b228;
    ram_cell[    8914] = 32'hbb307e90;
    ram_cell[    8915] = 32'hfbea23b0;
    ram_cell[    8916] = 32'h2c19f1aa;
    ram_cell[    8917] = 32'h5149dda6;
    ram_cell[    8918] = 32'h45cfd61d;
    ram_cell[    8919] = 32'h8cedf638;
    ram_cell[    8920] = 32'hdcbdc6d4;
    ram_cell[    8921] = 32'hbe51536e;
    ram_cell[    8922] = 32'ha938bff6;
    ram_cell[    8923] = 32'ha92e39d4;
    ram_cell[    8924] = 32'heedc28a8;
    ram_cell[    8925] = 32'h4d258a45;
    ram_cell[    8926] = 32'hf170929b;
    ram_cell[    8927] = 32'h6323349f;
    ram_cell[    8928] = 32'h9a7bd0a9;
    ram_cell[    8929] = 32'h8ecf35fc;
    ram_cell[    8930] = 32'h21c7b2b5;
    ram_cell[    8931] = 32'hc981f961;
    ram_cell[    8932] = 32'h6f10cb51;
    ram_cell[    8933] = 32'hff89ef57;
    ram_cell[    8934] = 32'hc287ad49;
    ram_cell[    8935] = 32'hf6b121a4;
    ram_cell[    8936] = 32'h06f52cb5;
    ram_cell[    8937] = 32'h978cf471;
    ram_cell[    8938] = 32'h8fe20a83;
    ram_cell[    8939] = 32'h86335c0b;
    ram_cell[    8940] = 32'he9bbed5b;
    ram_cell[    8941] = 32'h41ac11ce;
    ram_cell[    8942] = 32'ha2075d23;
    ram_cell[    8943] = 32'he0a12790;
    ram_cell[    8944] = 32'h6b504099;
    ram_cell[    8945] = 32'ha79deac9;
    ram_cell[    8946] = 32'h25e247d6;
    ram_cell[    8947] = 32'h4cbe015a;
    ram_cell[    8948] = 32'hdfb4a7ae;
    ram_cell[    8949] = 32'h361e3cf9;
    ram_cell[    8950] = 32'hd322cd13;
    ram_cell[    8951] = 32'h40cda42b;
    ram_cell[    8952] = 32'h30ae4e49;
    ram_cell[    8953] = 32'hc0ff68d6;
    ram_cell[    8954] = 32'h5cf9efbc;
    ram_cell[    8955] = 32'h80644727;
    ram_cell[    8956] = 32'h661f8246;
    ram_cell[    8957] = 32'hed2bb60d;
    ram_cell[    8958] = 32'h64e82a84;
    ram_cell[    8959] = 32'h96f0323b;
    ram_cell[    8960] = 32'he60639fd;
    ram_cell[    8961] = 32'h7a8e9c4c;
    ram_cell[    8962] = 32'hc518e54f;
    ram_cell[    8963] = 32'hb1593441;
    ram_cell[    8964] = 32'h6c1ff894;
    ram_cell[    8965] = 32'hcfb14206;
    ram_cell[    8966] = 32'hd38640f6;
    ram_cell[    8967] = 32'h835821d6;
    ram_cell[    8968] = 32'hea1a759e;
    ram_cell[    8969] = 32'h56f73dca;
    ram_cell[    8970] = 32'h73c53738;
    ram_cell[    8971] = 32'h41a4bd68;
    ram_cell[    8972] = 32'he854b53d;
    ram_cell[    8973] = 32'h1c6a965e;
    ram_cell[    8974] = 32'h049e1606;
    ram_cell[    8975] = 32'ha4328315;
    ram_cell[    8976] = 32'hbe50532a;
    ram_cell[    8977] = 32'hff191265;
    ram_cell[    8978] = 32'h74662746;
    ram_cell[    8979] = 32'h7c45882c;
    ram_cell[    8980] = 32'h32cc79be;
    ram_cell[    8981] = 32'h4796fdca;
    ram_cell[    8982] = 32'hf42ed56e;
    ram_cell[    8983] = 32'h2f962787;
    ram_cell[    8984] = 32'hb3f712b9;
    ram_cell[    8985] = 32'h72200898;
    ram_cell[    8986] = 32'hc175c3be;
    ram_cell[    8987] = 32'he352808f;
    ram_cell[    8988] = 32'h461be654;
    ram_cell[    8989] = 32'h04538574;
    ram_cell[    8990] = 32'h955b4450;
    ram_cell[    8991] = 32'h4ce2d112;
    ram_cell[    8992] = 32'h4ea06311;
    ram_cell[    8993] = 32'h293ba869;
    ram_cell[    8994] = 32'h0685a9b3;
    ram_cell[    8995] = 32'h6d4a1959;
    ram_cell[    8996] = 32'h0ed8255f;
    ram_cell[    8997] = 32'he6490b11;
    ram_cell[    8998] = 32'h7765d3f9;
    ram_cell[    8999] = 32'h99be7948;
    ram_cell[    9000] = 32'hf98dc138;
    ram_cell[    9001] = 32'hc0e161b5;
    ram_cell[    9002] = 32'h3ceb4bc7;
    ram_cell[    9003] = 32'ha3fa8ba4;
    ram_cell[    9004] = 32'h84858fa6;
    ram_cell[    9005] = 32'h9f73594a;
    ram_cell[    9006] = 32'haaf4ce08;
    ram_cell[    9007] = 32'hc15fb035;
    ram_cell[    9008] = 32'h6b06cf43;
    ram_cell[    9009] = 32'hf8c70c67;
    ram_cell[    9010] = 32'he5bb599d;
    ram_cell[    9011] = 32'h102d9a25;
    ram_cell[    9012] = 32'h022d3a89;
    ram_cell[    9013] = 32'h1777482a;
    ram_cell[    9014] = 32'h9bef6499;
    ram_cell[    9015] = 32'h9c8a2587;
    ram_cell[    9016] = 32'h757f47f4;
    ram_cell[    9017] = 32'h2f67c9c4;
    ram_cell[    9018] = 32'h7815c0a8;
    ram_cell[    9019] = 32'h65b0266e;
    ram_cell[    9020] = 32'hde437918;
    ram_cell[    9021] = 32'h75af8d5d;
    ram_cell[    9022] = 32'h650fe002;
    ram_cell[    9023] = 32'h20ff0151;
    ram_cell[    9024] = 32'h00bd39f3;
    ram_cell[    9025] = 32'h6cd9e62c;
    ram_cell[    9026] = 32'h7c4aaf4f;
    ram_cell[    9027] = 32'hb9133671;
    ram_cell[    9028] = 32'h09c987b1;
    ram_cell[    9029] = 32'hff259651;
    ram_cell[    9030] = 32'h4b2625e3;
    ram_cell[    9031] = 32'h2559efaf;
    ram_cell[    9032] = 32'h8a375924;
    ram_cell[    9033] = 32'hf5a8ea22;
    ram_cell[    9034] = 32'h046b13a9;
    ram_cell[    9035] = 32'h84e6b503;
    ram_cell[    9036] = 32'h978cef2f;
    ram_cell[    9037] = 32'h54a8aaed;
    ram_cell[    9038] = 32'he24dcbe4;
    ram_cell[    9039] = 32'he56885c1;
    ram_cell[    9040] = 32'h414f43c2;
    ram_cell[    9041] = 32'h7363c286;
    ram_cell[    9042] = 32'h1d4c1648;
    ram_cell[    9043] = 32'h5760f06a;
    ram_cell[    9044] = 32'h560dcb53;
    ram_cell[    9045] = 32'hac8a3874;
    ram_cell[    9046] = 32'h5a26faa2;
    ram_cell[    9047] = 32'hb68607aa;
    ram_cell[    9048] = 32'h7ba18895;
    ram_cell[    9049] = 32'h2772bcd9;
    ram_cell[    9050] = 32'h316d6096;
    ram_cell[    9051] = 32'h1f1eac97;
    ram_cell[    9052] = 32'h7ca5cef6;
    ram_cell[    9053] = 32'h40eb6998;
    ram_cell[    9054] = 32'h626dd050;
    ram_cell[    9055] = 32'h59f308b1;
    ram_cell[    9056] = 32'h5c0acee0;
    ram_cell[    9057] = 32'hcf3fd778;
    ram_cell[    9058] = 32'hc3840cc1;
    ram_cell[    9059] = 32'h41bb824f;
    ram_cell[    9060] = 32'h0e72d1d6;
    ram_cell[    9061] = 32'haf790dd8;
    ram_cell[    9062] = 32'h94655d8a;
    ram_cell[    9063] = 32'hae643af2;
    ram_cell[    9064] = 32'h054b5d5d;
    ram_cell[    9065] = 32'h663e7e01;
    ram_cell[    9066] = 32'h6eac8403;
    ram_cell[    9067] = 32'h3be9ce79;
    ram_cell[    9068] = 32'hc49dc303;
    ram_cell[    9069] = 32'h9520b7f1;
    ram_cell[    9070] = 32'h705a9765;
    ram_cell[    9071] = 32'hbc08043e;
    ram_cell[    9072] = 32'h14183a60;
    ram_cell[    9073] = 32'h8346fadf;
    ram_cell[    9074] = 32'hb3f82cb6;
    ram_cell[    9075] = 32'h3f507e0c;
    ram_cell[    9076] = 32'h8d982d49;
    ram_cell[    9077] = 32'hf04d8014;
    ram_cell[    9078] = 32'hc624718e;
    ram_cell[    9079] = 32'h3fe3a443;
    ram_cell[    9080] = 32'h460c6ced;
    ram_cell[    9081] = 32'h56db47db;
    ram_cell[    9082] = 32'h629317f2;
    ram_cell[    9083] = 32'h180fe219;
    ram_cell[    9084] = 32'h58e2d3ef;
    ram_cell[    9085] = 32'h04493cb4;
    ram_cell[    9086] = 32'hdfe581d2;
    ram_cell[    9087] = 32'hd9e2ff52;
    ram_cell[    9088] = 32'h62beb887;
    ram_cell[    9089] = 32'h3872cc05;
    ram_cell[    9090] = 32'ha8d0da5c;
    ram_cell[    9091] = 32'h5d3ee03f;
    ram_cell[    9092] = 32'ha8900a07;
    ram_cell[    9093] = 32'hf811bd9f;
    ram_cell[    9094] = 32'h0352a9f3;
    ram_cell[    9095] = 32'h12375d75;
    ram_cell[    9096] = 32'h35ee0a9b;
    ram_cell[    9097] = 32'h2b9ea833;
    ram_cell[    9098] = 32'hcaa9a288;
    ram_cell[    9099] = 32'h64184e3e;
    ram_cell[    9100] = 32'hd9a81a4d;
    ram_cell[    9101] = 32'h9f67e392;
    ram_cell[    9102] = 32'hba2acdf2;
    ram_cell[    9103] = 32'h18a8dbed;
    ram_cell[    9104] = 32'h70556106;
    ram_cell[    9105] = 32'h3f177df2;
    ram_cell[    9106] = 32'h2e21aae1;
    ram_cell[    9107] = 32'h4ee026b3;
    ram_cell[    9108] = 32'h2d63fc9d;
    ram_cell[    9109] = 32'h2cf6a493;
    ram_cell[    9110] = 32'h7a54ed98;
    ram_cell[    9111] = 32'h871f0f83;
    ram_cell[    9112] = 32'heab905a8;
    ram_cell[    9113] = 32'h7c51a426;
    ram_cell[    9114] = 32'h107a5e46;
    ram_cell[    9115] = 32'hf2795655;
    ram_cell[    9116] = 32'h0d15f279;
    ram_cell[    9117] = 32'h6926bc1d;
    ram_cell[    9118] = 32'h74ee0dd3;
    ram_cell[    9119] = 32'h96f9771f;
    ram_cell[    9120] = 32'h0b8d4b51;
    ram_cell[    9121] = 32'hb733efb6;
    ram_cell[    9122] = 32'hee13f7d6;
    ram_cell[    9123] = 32'h72f48146;
    ram_cell[    9124] = 32'hafbbf1d0;
    ram_cell[    9125] = 32'h9009eb82;
    ram_cell[    9126] = 32'h9ff8bc33;
    ram_cell[    9127] = 32'h99e30824;
    ram_cell[    9128] = 32'ha6f3f731;
    ram_cell[    9129] = 32'hae17f233;
    ram_cell[    9130] = 32'hc6b8e3a9;
    ram_cell[    9131] = 32'he66d4ce4;
    ram_cell[    9132] = 32'h7b3ba6ff;
    ram_cell[    9133] = 32'hb0d3f1ca;
    ram_cell[    9134] = 32'hbb5a9acf;
    ram_cell[    9135] = 32'h6d1c9065;
    ram_cell[    9136] = 32'hfc864b6f;
    ram_cell[    9137] = 32'h3b2705d5;
    ram_cell[    9138] = 32'h8d74d184;
    ram_cell[    9139] = 32'h4217731e;
    ram_cell[    9140] = 32'hc8cae34e;
    ram_cell[    9141] = 32'h2d229e1a;
    ram_cell[    9142] = 32'h48656db0;
    ram_cell[    9143] = 32'h87ae821f;
    ram_cell[    9144] = 32'h72349c59;
    ram_cell[    9145] = 32'hdeaba4e0;
    ram_cell[    9146] = 32'h2ac3c524;
    ram_cell[    9147] = 32'h3b7150b9;
    ram_cell[    9148] = 32'had301909;
    ram_cell[    9149] = 32'h3507d508;
    ram_cell[    9150] = 32'h2d2b7363;
    ram_cell[    9151] = 32'h24c9b43e;
    ram_cell[    9152] = 32'h63205e2c;
    ram_cell[    9153] = 32'ha1653934;
    ram_cell[    9154] = 32'h313f2bc2;
    ram_cell[    9155] = 32'hc7e14869;
    ram_cell[    9156] = 32'he7ae074e;
    ram_cell[    9157] = 32'hd99ebf56;
    ram_cell[    9158] = 32'h93d509d2;
    ram_cell[    9159] = 32'h67c364d1;
    ram_cell[    9160] = 32'he98d9c08;
    ram_cell[    9161] = 32'hc2621274;
    ram_cell[    9162] = 32'h2fab5150;
    ram_cell[    9163] = 32'h0a2e4a33;
    ram_cell[    9164] = 32'ha2fac8f1;
    ram_cell[    9165] = 32'hf852f739;
    ram_cell[    9166] = 32'hecd6d214;
    ram_cell[    9167] = 32'h9d76ff0f;
    ram_cell[    9168] = 32'hb9b3e73f;
    ram_cell[    9169] = 32'hf74d752a;
    ram_cell[    9170] = 32'h4c600928;
    ram_cell[    9171] = 32'h322cea52;
    ram_cell[    9172] = 32'h53267b08;
    ram_cell[    9173] = 32'h355b9f3e;
    ram_cell[    9174] = 32'h14d4c8c8;
    ram_cell[    9175] = 32'h2eaa2348;
    ram_cell[    9176] = 32'hea67d658;
    ram_cell[    9177] = 32'hedc7f2bf;
    ram_cell[    9178] = 32'hc8599b83;
    ram_cell[    9179] = 32'h1bb0a51d;
    ram_cell[    9180] = 32'h8d791e74;
    ram_cell[    9181] = 32'h04d544f7;
    ram_cell[    9182] = 32'h0f066399;
    ram_cell[    9183] = 32'h5027e2e9;
    ram_cell[    9184] = 32'hec79ab68;
    ram_cell[    9185] = 32'hc32535f0;
    ram_cell[    9186] = 32'h660c2025;
    ram_cell[    9187] = 32'hff83c6c8;
    ram_cell[    9188] = 32'he377fc71;
    ram_cell[    9189] = 32'h33a450f8;
    ram_cell[    9190] = 32'hdc3d5b23;
    ram_cell[    9191] = 32'hd2acfad8;
    ram_cell[    9192] = 32'hc2fde593;
    ram_cell[    9193] = 32'he1489b39;
    ram_cell[    9194] = 32'hfda6164b;
    ram_cell[    9195] = 32'h411ac9c9;
    ram_cell[    9196] = 32'h99521570;
    ram_cell[    9197] = 32'h76867328;
    ram_cell[    9198] = 32'h7649a4bb;
    ram_cell[    9199] = 32'h2c936e18;
    ram_cell[    9200] = 32'h7e29dedd;
    ram_cell[    9201] = 32'hcdfa3cfb;
    ram_cell[    9202] = 32'h5ffa49df;
    ram_cell[    9203] = 32'h2aab273a;
    ram_cell[    9204] = 32'h894677c7;
    ram_cell[    9205] = 32'h6836a71a;
    ram_cell[    9206] = 32'h533d8a42;
    ram_cell[    9207] = 32'h76b48c2c;
    ram_cell[    9208] = 32'h99786fcb;
    ram_cell[    9209] = 32'hc5e0fcef;
    ram_cell[    9210] = 32'h9a010846;
    ram_cell[    9211] = 32'h53d478b7;
    ram_cell[    9212] = 32'h45a9b0f5;
    ram_cell[    9213] = 32'h00dd5a47;
    ram_cell[    9214] = 32'h41b47e9d;
    ram_cell[    9215] = 32'h9394da73;
    ram_cell[    9216] = 32'hafac7ad2;
    ram_cell[    9217] = 32'h10e5ab8b;
    ram_cell[    9218] = 32'hbd7d9662;
    ram_cell[    9219] = 32'hc2cf1575;
    ram_cell[    9220] = 32'h229fb200;
    ram_cell[    9221] = 32'h0737386e;
    ram_cell[    9222] = 32'ha436b567;
    ram_cell[    9223] = 32'h9d7bb3b7;
    ram_cell[    9224] = 32'hd1929a8b;
    ram_cell[    9225] = 32'hf0ff228a;
    ram_cell[    9226] = 32'hc611d8cc;
    ram_cell[    9227] = 32'hf7160e76;
    ram_cell[    9228] = 32'h254a2c32;
    ram_cell[    9229] = 32'hc84c547f;
    ram_cell[    9230] = 32'h4b42399d;
    ram_cell[    9231] = 32'h436b228e;
    ram_cell[    9232] = 32'hbe78c662;
    ram_cell[    9233] = 32'h342c83c1;
    ram_cell[    9234] = 32'he6396891;
    ram_cell[    9235] = 32'h957c78eb;
    ram_cell[    9236] = 32'h820ef906;
    ram_cell[    9237] = 32'h126f1be0;
    ram_cell[    9238] = 32'hea319517;
    ram_cell[    9239] = 32'h6a67a6ac;
    ram_cell[    9240] = 32'ha08049ee;
    ram_cell[    9241] = 32'hc89acbc1;
    ram_cell[    9242] = 32'h16fef320;
    ram_cell[    9243] = 32'h040c9333;
    ram_cell[    9244] = 32'h5dde7dfa;
    ram_cell[    9245] = 32'ha88689c3;
    ram_cell[    9246] = 32'h8b18d062;
    ram_cell[    9247] = 32'h8eb2061c;
    ram_cell[    9248] = 32'h1b815eb1;
    ram_cell[    9249] = 32'ha6d0a478;
    ram_cell[    9250] = 32'h34479841;
    ram_cell[    9251] = 32'h916cc222;
    ram_cell[    9252] = 32'hfd56a6be;
    ram_cell[    9253] = 32'ha8ec5dc8;
    ram_cell[    9254] = 32'h58001bc7;
    ram_cell[    9255] = 32'hf259ebc5;
    ram_cell[    9256] = 32'h98b7e629;
    ram_cell[    9257] = 32'hf0454176;
    ram_cell[    9258] = 32'hd70b5810;
    ram_cell[    9259] = 32'h147c3f9a;
    ram_cell[    9260] = 32'h574aab13;
    ram_cell[    9261] = 32'hd7bab2e1;
    ram_cell[    9262] = 32'hd7260375;
    ram_cell[    9263] = 32'h745e06f9;
    ram_cell[    9264] = 32'he37e381c;
    ram_cell[    9265] = 32'h94679438;
    ram_cell[    9266] = 32'h8de9133e;
    ram_cell[    9267] = 32'hd6b0e1b0;
    ram_cell[    9268] = 32'h2fab7ffa;
    ram_cell[    9269] = 32'h6924ec43;
    ram_cell[    9270] = 32'hc2a40a60;
    ram_cell[    9271] = 32'h9105b608;
    ram_cell[    9272] = 32'hdfad8359;
    ram_cell[    9273] = 32'h7e1d4a48;
    ram_cell[    9274] = 32'h2f526752;
    ram_cell[    9275] = 32'hf9d54eb0;
    ram_cell[    9276] = 32'h165188c0;
    ram_cell[    9277] = 32'hf1dcac90;
    ram_cell[    9278] = 32'h63a91524;
    ram_cell[    9279] = 32'hdf82d57d;
    ram_cell[    9280] = 32'h8c070828;
    ram_cell[    9281] = 32'h5015c088;
    ram_cell[    9282] = 32'hc96ccec1;
    ram_cell[    9283] = 32'hf6fd7ec2;
    ram_cell[    9284] = 32'hefa3269b;
    ram_cell[    9285] = 32'h94738926;
    ram_cell[    9286] = 32'h761daa54;
    ram_cell[    9287] = 32'h759d992b;
    ram_cell[    9288] = 32'hd1fefc62;
    ram_cell[    9289] = 32'h182ca355;
    ram_cell[    9290] = 32'hef5794b7;
    ram_cell[    9291] = 32'h130ac3b1;
    ram_cell[    9292] = 32'h4fbc8406;
    ram_cell[    9293] = 32'h56115b34;
    ram_cell[    9294] = 32'hfacc10ae;
    ram_cell[    9295] = 32'ha34b8114;
    ram_cell[    9296] = 32'h30bfe388;
    ram_cell[    9297] = 32'hcfa58148;
    ram_cell[    9298] = 32'he89b73b3;
    ram_cell[    9299] = 32'ha12f2e0a;
    ram_cell[    9300] = 32'h2353181f;
    ram_cell[    9301] = 32'h2d373eed;
    ram_cell[    9302] = 32'h32890471;
    ram_cell[    9303] = 32'ha9e10b69;
    ram_cell[    9304] = 32'h669c19b0;
    ram_cell[    9305] = 32'he0ba8946;
    ram_cell[    9306] = 32'h62880c6c;
    ram_cell[    9307] = 32'h290ac810;
    ram_cell[    9308] = 32'hd6909089;
    ram_cell[    9309] = 32'hcffc9763;
    ram_cell[    9310] = 32'h0df4a22b;
    ram_cell[    9311] = 32'h17a1ee66;
    ram_cell[    9312] = 32'hddfc08c2;
    ram_cell[    9313] = 32'h3fa9f2e7;
    ram_cell[    9314] = 32'hc2020e72;
    ram_cell[    9315] = 32'hd86f9ccb;
    ram_cell[    9316] = 32'h708f996b;
    ram_cell[    9317] = 32'h0143b91d;
    ram_cell[    9318] = 32'hca25737e;
    ram_cell[    9319] = 32'hc425378a;
    ram_cell[    9320] = 32'ha7f301df;
    ram_cell[    9321] = 32'h1a99c2fe;
    ram_cell[    9322] = 32'ha981d7ce;
    ram_cell[    9323] = 32'hb24794ed;
    ram_cell[    9324] = 32'h6a18b096;
    ram_cell[    9325] = 32'he3f471c8;
    ram_cell[    9326] = 32'hf063ac46;
    ram_cell[    9327] = 32'h55cf3db0;
    ram_cell[    9328] = 32'hafde8890;
    ram_cell[    9329] = 32'h4cf0ab07;
    ram_cell[    9330] = 32'haa48b29d;
    ram_cell[    9331] = 32'hf3a0b47e;
    ram_cell[    9332] = 32'ha0492643;
    ram_cell[    9333] = 32'h61a89f1c;
    ram_cell[    9334] = 32'h6690d9f7;
    ram_cell[    9335] = 32'h109f91d3;
    ram_cell[    9336] = 32'h136844aa;
    ram_cell[    9337] = 32'h9334b349;
    ram_cell[    9338] = 32'h084c955f;
    ram_cell[    9339] = 32'hc64cd07f;
    ram_cell[    9340] = 32'h96024b2a;
    ram_cell[    9341] = 32'h0774cace;
    ram_cell[    9342] = 32'hb8278d9a;
    ram_cell[    9343] = 32'he640ed26;
    ram_cell[    9344] = 32'hfea8bdd6;
    ram_cell[    9345] = 32'h962f244f;
    ram_cell[    9346] = 32'h86ba4d25;
    ram_cell[    9347] = 32'hcd71efb1;
    ram_cell[    9348] = 32'hcebf3a9b;
    ram_cell[    9349] = 32'h5372d144;
    ram_cell[    9350] = 32'h86d12650;
    ram_cell[    9351] = 32'h1257ea06;
    ram_cell[    9352] = 32'h6e4a3285;
    ram_cell[    9353] = 32'h593c2768;
    ram_cell[    9354] = 32'h34aa7ab1;
    ram_cell[    9355] = 32'h3576caba;
    ram_cell[    9356] = 32'he6af1fef;
    ram_cell[    9357] = 32'h90416a6f;
    ram_cell[    9358] = 32'h8a4ce11d;
    ram_cell[    9359] = 32'h11d3c6a4;
    ram_cell[    9360] = 32'h3d864092;
    ram_cell[    9361] = 32'h7e20f5a1;
    ram_cell[    9362] = 32'h8a809e1a;
    ram_cell[    9363] = 32'h0c99d615;
    ram_cell[    9364] = 32'hd6412a91;
    ram_cell[    9365] = 32'h1c5d748e;
    ram_cell[    9366] = 32'h8714933b;
    ram_cell[    9367] = 32'h5a0f15b5;
    ram_cell[    9368] = 32'h0a9318ef;
    ram_cell[    9369] = 32'h45cab000;
    ram_cell[    9370] = 32'h754029a0;
    ram_cell[    9371] = 32'h4fafd6a3;
    ram_cell[    9372] = 32'hbfb8c03d;
    ram_cell[    9373] = 32'h08e3d215;
    ram_cell[    9374] = 32'h0897d722;
    ram_cell[    9375] = 32'h27d41e12;
    ram_cell[    9376] = 32'hecf00f8d;
    ram_cell[    9377] = 32'h50fda83c;
    ram_cell[    9378] = 32'h68d577c2;
    ram_cell[    9379] = 32'h5bd687a1;
    ram_cell[    9380] = 32'h03d712b0;
    ram_cell[    9381] = 32'h883b1ede;
    ram_cell[    9382] = 32'h4fc6b2ff;
    ram_cell[    9383] = 32'hc128de12;
    ram_cell[    9384] = 32'h84787e70;
    ram_cell[    9385] = 32'h8548e72c;
    ram_cell[    9386] = 32'he56ca574;
    ram_cell[    9387] = 32'h537338c9;
    ram_cell[    9388] = 32'h77f5857d;
    ram_cell[    9389] = 32'hedae31f9;
    ram_cell[    9390] = 32'h08651045;
    ram_cell[    9391] = 32'hf622c35e;
    ram_cell[    9392] = 32'hdc67dc7d;
    ram_cell[    9393] = 32'h6cf42598;
    ram_cell[    9394] = 32'h93158b88;
    ram_cell[    9395] = 32'h6ff8a502;
    ram_cell[    9396] = 32'hacdc8162;
    ram_cell[    9397] = 32'hc6cb32f7;
    ram_cell[    9398] = 32'h981e4a7c;
    ram_cell[    9399] = 32'h5e93c516;
    ram_cell[    9400] = 32'h1e6bd30d;
    ram_cell[    9401] = 32'hef89aeb4;
    ram_cell[    9402] = 32'h1f373090;
    ram_cell[    9403] = 32'hac959a88;
    ram_cell[    9404] = 32'h6bb05bcb;
    ram_cell[    9405] = 32'h935cf1e8;
    ram_cell[    9406] = 32'he8632088;
    ram_cell[    9407] = 32'hdb563afb;
    ram_cell[    9408] = 32'h8ef6c375;
    ram_cell[    9409] = 32'he0790352;
    ram_cell[    9410] = 32'ha1c7a3b8;
    ram_cell[    9411] = 32'h72cb3a79;
    ram_cell[    9412] = 32'h0e48c70f;
    ram_cell[    9413] = 32'hbe7e50b3;
    ram_cell[    9414] = 32'h8f544387;
    ram_cell[    9415] = 32'hc5660869;
    ram_cell[    9416] = 32'h0dcc8135;
    ram_cell[    9417] = 32'h593b1c41;
    ram_cell[    9418] = 32'h0108d0d9;
    ram_cell[    9419] = 32'hbcf29473;
    ram_cell[    9420] = 32'h166a0549;
    ram_cell[    9421] = 32'h724eab45;
    ram_cell[    9422] = 32'he88596d2;
    ram_cell[    9423] = 32'ha2ee76aa;
    ram_cell[    9424] = 32'hd1b8f861;
    ram_cell[    9425] = 32'h4f310e5e;
    ram_cell[    9426] = 32'h1111bcad;
    ram_cell[    9427] = 32'h054bc534;
    ram_cell[    9428] = 32'hc67b9b02;
    ram_cell[    9429] = 32'h226eccaf;
    ram_cell[    9430] = 32'hc26cfe67;
    ram_cell[    9431] = 32'he73216fc;
    ram_cell[    9432] = 32'h9611a9a9;
    ram_cell[    9433] = 32'h8bfa16c2;
    ram_cell[    9434] = 32'hd3de5f3e;
    ram_cell[    9435] = 32'h021c8973;
    ram_cell[    9436] = 32'h12e483db;
    ram_cell[    9437] = 32'he522e693;
    ram_cell[    9438] = 32'hd94f4fa1;
    ram_cell[    9439] = 32'hcae3ec78;
    ram_cell[    9440] = 32'h2ea527b0;
    ram_cell[    9441] = 32'h13319e55;
    ram_cell[    9442] = 32'he35fef17;
    ram_cell[    9443] = 32'hc061371d;
    ram_cell[    9444] = 32'hb155c619;
    ram_cell[    9445] = 32'h5222a004;
    ram_cell[    9446] = 32'h54b7d76c;
    ram_cell[    9447] = 32'h7a38b23e;
    ram_cell[    9448] = 32'h4efab43d;
    ram_cell[    9449] = 32'h163d5146;
    ram_cell[    9450] = 32'h76f37e7e;
    ram_cell[    9451] = 32'h77530641;
    ram_cell[    9452] = 32'h02dd6577;
    ram_cell[    9453] = 32'h671a311f;
    ram_cell[    9454] = 32'hcced2ec2;
    ram_cell[    9455] = 32'h002ad8e3;
    ram_cell[    9456] = 32'hc47cbdac;
    ram_cell[    9457] = 32'h5fa6e8a5;
    ram_cell[    9458] = 32'h9219bd55;
    ram_cell[    9459] = 32'h8cef04ed;
    ram_cell[    9460] = 32'hc3186761;
    ram_cell[    9461] = 32'he13ddd6c;
    ram_cell[    9462] = 32'hb4c3d22e;
    ram_cell[    9463] = 32'h68dfc4ac;
    ram_cell[    9464] = 32'h4e3d2729;
    ram_cell[    9465] = 32'hced57b46;
    ram_cell[    9466] = 32'hd3489388;
    ram_cell[    9467] = 32'h02da1e32;
    ram_cell[    9468] = 32'haa88a3eb;
    ram_cell[    9469] = 32'h5e1630c3;
    ram_cell[    9470] = 32'hfebc89f8;
    ram_cell[    9471] = 32'ha9317821;
    ram_cell[    9472] = 32'h9448137c;
    ram_cell[    9473] = 32'h2cbf7732;
    ram_cell[    9474] = 32'h419e3878;
    ram_cell[    9475] = 32'hb7ace417;
    ram_cell[    9476] = 32'h5692716a;
    ram_cell[    9477] = 32'h31423dda;
    ram_cell[    9478] = 32'h644944ec;
    ram_cell[    9479] = 32'h44872179;
    ram_cell[    9480] = 32'hda4a6a3f;
    ram_cell[    9481] = 32'h32aa6cdc;
    ram_cell[    9482] = 32'h2025652d;
    ram_cell[    9483] = 32'h4f6b07a3;
    ram_cell[    9484] = 32'had9afa72;
    ram_cell[    9485] = 32'h89919670;
    ram_cell[    9486] = 32'hc445c3e4;
    ram_cell[    9487] = 32'h3b07dd5e;
    ram_cell[    9488] = 32'h135558d8;
    ram_cell[    9489] = 32'h03d23812;
    ram_cell[    9490] = 32'h55424bd0;
    ram_cell[    9491] = 32'haf42788e;
    ram_cell[    9492] = 32'h2e542c66;
    ram_cell[    9493] = 32'h0654aa43;
    ram_cell[    9494] = 32'hb7f9dba7;
    ram_cell[    9495] = 32'h21c7cb3c;
    ram_cell[    9496] = 32'h3f38c59c;
    ram_cell[    9497] = 32'hc985cd52;
    ram_cell[    9498] = 32'h04904fd4;
    ram_cell[    9499] = 32'h82531b99;
    ram_cell[    9500] = 32'h7c2a9e09;
    ram_cell[    9501] = 32'h0a1e9a45;
    ram_cell[    9502] = 32'h48f97dd7;
    ram_cell[    9503] = 32'hfc720658;
    ram_cell[    9504] = 32'h8fa6fa39;
    ram_cell[    9505] = 32'h76e297b7;
    ram_cell[    9506] = 32'h326a994c;
    ram_cell[    9507] = 32'hdb46772c;
    ram_cell[    9508] = 32'h4043975d;
    ram_cell[    9509] = 32'h26fd2457;
    ram_cell[    9510] = 32'h188602fa;
    ram_cell[    9511] = 32'h158986ea;
    ram_cell[    9512] = 32'h10ca8fc2;
    ram_cell[    9513] = 32'h5dce40db;
    ram_cell[    9514] = 32'hcc280531;
    ram_cell[    9515] = 32'h8fa73e8c;
    ram_cell[    9516] = 32'h9b5b6470;
    ram_cell[    9517] = 32'h8d0586b2;
    ram_cell[    9518] = 32'haaad98b3;
    ram_cell[    9519] = 32'heb4b9acd;
    ram_cell[    9520] = 32'h77135729;
    ram_cell[    9521] = 32'hc2553900;
    ram_cell[    9522] = 32'h0ffde5a5;
    ram_cell[    9523] = 32'h7cb4bf1a;
    ram_cell[    9524] = 32'hf4740566;
    ram_cell[    9525] = 32'h22894bab;
    ram_cell[    9526] = 32'h002dfcd6;
    ram_cell[    9527] = 32'h3a63b55e;
    ram_cell[    9528] = 32'h7bea00c2;
    ram_cell[    9529] = 32'hf38b0482;
    ram_cell[    9530] = 32'h6398d729;
    ram_cell[    9531] = 32'h74ae95e6;
    ram_cell[    9532] = 32'hdc6b7927;
    ram_cell[    9533] = 32'hbbed4f05;
    ram_cell[    9534] = 32'hdb35a82f;
    ram_cell[    9535] = 32'h754d8017;
    ram_cell[    9536] = 32'h533e21d9;
    ram_cell[    9537] = 32'h1ca6492d;
    ram_cell[    9538] = 32'h43d99302;
    ram_cell[    9539] = 32'he39645e2;
    ram_cell[    9540] = 32'hf2ca66f5;
    ram_cell[    9541] = 32'h5160ed33;
    ram_cell[    9542] = 32'hbc66c632;
    ram_cell[    9543] = 32'h5f96f9cf;
    ram_cell[    9544] = 32'h876ac7db;
    ram_cell[    9545] = 32'h8c257f87;
    ram_cell[    9546] = 32'hb28949a7;
    ram_cell[    9547] = 32'ha2736ed8;
    ram_cell[    9548] = 32'h58116318;
    ram_cell[    9549] = 32'h1c1831b1;
    ram_cell[    9550] = 32'heaffb0ac;
    ram_cell[    9551] = 32'h99063ad8;
    ram_cell[    9552] = 32'h4fa05c42;
    ram_cell[    9553] = 32'h7c51feb1;
    ram_cell[    9554] = 32'h416e5546;
    ram_cell[    9555] = 32'h2a2201c7;
    ram_cell[    9556] = 32'h4e566604;
    ram_cell[    9557] = 32'h9ba8ffe4;
    ram_cell[    9558] = 32'h361e6d67;
    ram_cell[    9559] = 32'h33cec80a;
    ram_cell[    9560] = 32'hb6a87f9e;
    ram_cell[    9561] = 32'hb845c8f6;
    ram_cell[    9562] = 32'hc5616c2e;
    ram_cell[    9563] = 32'h7c09cc4a;
    ram_cell[    9564] = 32'h716e93bb;
    ram_cell[    9565] = 32'hf8d59f98;
    ram_cell[    9566] = 32'h0f7d4e62;
    ram_cell[    9567] = 32'h7894f1c3;
    ram_cell[    9568] = 32'hd437b86a;
    ram_cell[    9569] = 32'h0655a144;
    ram_cell[    9570] = 32'h1965d93c;
    ram_cell[    9571] = 32'h1dca7d7e;
    ram_cell[    9572] = 32'h44a1536d;
    ram_cell[    9573] = 32'hd5f48964;
    ram_cell[    9574] = 32'h83b9b637;
    ram_cell[    9575] = 32'h4383e976;
    ram_cell[    9576] = 32'h40b6169b;
    ram_cell[    9577] = 32'hb4133599;
    ram_cell[    9578] = 32'hc89ac00d;
    ram_cell[    9579] = 32'h8725cb77;
    ram_cell[    9580] = 32'h787ad00d;
    ram_cell[    9581] = 32'he7c23ebe;
    ram_cell[    9582] = 32'ha5852913;
    ram_cell[    9583] = 32'h99952bf6;
    ram_cell[    9584] = 32'hf9df5916;
    ram_cell[    9585] = 32'h1c4c9183;
    ram_cell[    9586] = 32'hfb0a25e6;
    ram_cell[    9587] = 32'h71989751;
    ram_cell[    9588] = 32'hd9c548a4;
    ram_cell[    9589] = 32'he1a1aa0b;
    ram_cell[    9590] = 32'hc79dc3c8;
    ram_cell[    9591] = 32'h68716891;
    ram_cell[    9592] = 32'hddf1cc3b;
    ram_cell[    9593] = 32'h0ae13dfc;
    ram_cell[    9594] = 32'hc04d2db9;
    ram_cell[    9595] = 32'hafc60f95;
    ram_cell[    9596] = 32'hf0d1fec7;
    ram_cell[    9597] = 32'he7abd429;
    ram_cell[    9598] = 32'hc6da2e98;
    ram_cell[    9599] = 32'h9fb38472;
    ram_cell[    9600] = 32'h270681b3;
    ram_cell[    9601] = 32'h7953386f;
    ram_cell[    9602] = 32'h84304641;
    ram_cell[    9603] = 32'hfbcfd3ab;
    ram_cell[    9604] = 32'h06345b69;
    ram_cell[    9605] = 32'h405be552;
    ram_cell[    9606] = 32'h6dc8d717;
    ram_cell[    9607] = 32'hde98bbb8;
    ram_cell[    9608] = 32'hb1266348;
    ram_cell[    9609] = 32'h3a68cdfa;
    ram_cell[    9610] = 32'h612006a0;
    ram_cell[    9611] = 32'h5f6834b8;
    ram_cell[    9612] = 32'hc5b9b570;
    ram_cell[    9613] = 32'hee7bd549;
    ram_cell[    9614] = 32'h3e3ff6e9;
    ram_cell[    9615] = 32'h203b70b1;
    ram_cell[    9616] = 32'ha7434c93;
    ram_cell[    9617] = 32'hcff48c40;
    ram_cell[    9618] = 32'h541d21ab;
    ram_cell[    9619] = 32'h756ea796;
    ram_cell[    9620] = 32'he2a2248f;
    ram_cell[    9621] = 32'h94253e48;
    ram_cell[    9622] = 32'hddbbe49f;
    ram_cell[    9623] = 32'h18bf6dc4;
    ram_cell[    9624] = 32'hc7c990cb;
    ram_cell[    9625] = 32'h23d46213;
    ram_cell[    9626] = 32'h89c1fb20;
    ram_cell[    9627] = 32'hd68e6118;
    ram_cell[    9628] = 32'h75b22af6;
    ram_cell[    9629] = 32'h25d19d88;
    ram_cell[    9630] = 32'h6a6fcb67;
    ram_cell[    9631] = 32'h8e788dbd;
    ram_cell[    9632] = 32'hc9b5fdfa;
    ram_cell[    9633] = 32'h4a3f8874;
    ram_cell[    9634] = 32'hec33ea28;
    ram_cell[    9635] = 32'h1e0da093;
    ram_cell[    9636] = 32'h647c4658;
    ram_cell[    9637] = 32'h4fc5bf22;
    ram_cell[    9638] = 32'h62d1758b;
    ram_cell[    9639] = 32'h615f43f0;
    ram_cell[    9640] = 32'h4e7afea9;
    ram_cell[    9641] = 32'hb3a095e8;
    ram_cell[    9642] = 32'hf2c715e6;
    ram_cell[    9643] = 32'heb1d794d;
    ram_cell[    9644] = 32'hee400b20;
    ram_cell[    9645] = 32'he6c0efe1;
    ram_cell[    9646] = 32'h7a4387ad;
    ram_cell[    9647] = 32'h6877d40f;
    ram_cell[    9648] = 32'hd0668498;
    ram_cell[    9649] = 32'h1583b5d4;
    ram_cell[    9650] = 32'h5389fd9f;
    ram_cell[    9651] = 32'hdbae4549;
    ram_cell[    9652] = 32'h04894825;
    ram_cell[    9653] = 32'h3d1559d0;
    ram_cell[    9654] = 32'he479b90c;
    ram_cell[    9655] = 32'h48abfee3;
    ram_cell[    9656] = 32'h5ba37eb3;
    ram_cell[    9657] = 32'h95f350a4;
    ram_cell[    9658] = 32'h0f046c0c;
    ram_cell[    9659] = 32'hf6a55fd1;
    ram_cell[    9660] = 32'hcac64ea3;
    ram_cell[    9661] = 32'h3b7c6e68;
    ram_cell[    9662] = 32'hd21dc492;
    ram_cell[    9663] = 32'h5546e388;
    ram_cell[    9664] = 32'h91f1d5d3;
    ram_cell[    9665] = 32'hb6af01af;
    ram_cell[    9666] = 32'h49ad2c49;
    ram_cell[    9667] = 32'h4bae75c5;
    ram_cell[    9668] = 32'h162144e4;
    ram_cell[    9669] = 32'hcc2b7fae;
    ram_cell[    9670] = 32'h52bb37e5;
    ram_cell[    9671] = 32'hbebadf7c;
    ram_cell[    9672] = 32'h758bbfd2;
    ram_cell[    9673] = 32'he4252ab0;
    ram_cell[    9674] = 32'hb191d779;
    ram_cell[    9675] = 32'h82196161;
    ram_cell[    9676] = 32'h175cd60d;
    ram_cell[    9677] = 32'h573455fc;
    ram_cell[    9678] = 32'hd3eafcd2;
    ram_cell[    9679] = 32'h09cfe75c;
    ram_cell[    9680] = 32'h20cb25d7;
    ram_cell[    9681] = 32'h1c78a1db;
    ram_cell[    9682] = 32'h2cbba526;
    ram_cell[    9683] = 32'h6487ba20;
    ram_cell[    9684] = 32'h4066c87c;
    ram_cell[    9685] = 32'hbc7b5077;
    ram_cell[    9686] = 32'h3aac323c;
    ram_cell[    9687] = 32'h7a1ed1ee;
    ram_cell[    9688] = 32'hb9cd9c7c;
    ram_cell[    9689] = 32'h4bed28f1;
    ram_cell[    9690] = 32'h1031e904;
    ram_cell[    9691] = 32'hb5ab4e48;
    ram_cell[    9692] = 32'hf658f0e5;
    ram_cell[    9693] = 32'h8eb9df4b;
    ram_cell[    9694] = 32'h0c186b15;
    ram_cell[    9695] = 32'h79f17f30;
    ram_cell[    9696] = 32'h5a1048c5;
    ram_cell[    9697] = 32'h714b13b1;
    ram_cell[    9698] = 32'h420e1d6a;
    ram_cell[    9699] = 32'h6f88a426;
    ram_cell[    9700] = 32'hae4f8f4d;
    ram_cell[    9701] = 32'h20c0aab7;
    ram_cell[    9702] = 32'h4a0c497a;
    ram_cell[    9703] = 32'h7c1e79a3;
    ram_cell[    9704] = 32'hae8fd2f0;
    ram_cell[    9705] = 32'hf52bfc09;
    ram_cell[    9706] = 32'h43f4c97b;
    ram_cell[    9707] = 32'h08d8df40;
    ram_cell[    9708] = 32'he22a2e54;
    ram_cell[    9709] = 32'hea45aff9;
    ram_cell[    9710] = 32'h52be250f;
    ram_cell[    9711] = 32'h23bafaf2;
    ram_cell[    9712] = 32'had0d4d30;
    ram_cell[    9713] = 32'hf35c4b4f;
    ram_cell[    9714] = 32'h4aa1359a;
    ram_cell[    9715] = 32'h6683979d;
    ram_cell[    9716] = 32'hd76b4835;
    ram_cell[    9717] = 32'hcf0d729a;
    ram_cell[    9718] = 32'h0d5d98c1;
    ram_cell[    9719] = 32'h28816bab;
    ram_cell[    9720] = 32'h5fb66e22;
    ram_cell[    9721] = 32'hf3536189;
    ram_cell[    9722] = 32'h8d9f7611;
    ram_cell[    9723] = 32'hb38069b4;
    ram_cell[    9724] = 32'ha7699127;
    ram_cell[    9725] = 32'he3c6685c;
    ram_cell[    9726] = 32'h0a5bb3b9;
    ram_cell[    9727] = 32'h9be18343;
    ram_cell[    9728] = 32'h4d0642bf;
    ram_cell[    9729] = 32'hed81ea92;
    ram_cell[    9730] = 32'hc8faf6a6;
    ram_cell[    9731] = 32'he51abdd6;
    ram_cell[    9732] = 32'hf5541d43;
    ram_cell[    9733] = 32'heed02711;
    ram_cell[    9734] = 32'h7c4720e9;
    ram_cell[    9735] = 32'h88c981eb;
    ram_cell[    9736] = 32'hf581a7c0;
    ram_cell[    9737] = 32'h7c8f0591;
    ram_cell[    9738] = 32'h8e5d19df;
    ram_cell[    9739] = 32'h00766f04;
    ram_cell[    9740] = 32'hc046b6d7;
    ram_cell[    9741] = 32'ha3d55995;
    ram_cell[    9742] = 32'h4863007a;
    ram_cell[    9743] = 32'h78c0460c;
    ram_cell[    9744] = 32'h90a7cee3;
    ram_cell[    9745] = 32'h1ed1e813;
    ram_cell[    9746] = 32'h9ebbd7ad;
    ram_cell[    9747] = 32'h4079f796;
    ram_cell[    9748] = 32'h314a503c;
    ram_cell[    9749] = 32'ha882b3d3;
    ram_cell[    9750] = 32'hccb603d7;
    ram_cell[    9751] = 32'h8747267c;
    ram_cell[    9752] = 32'hb66ea72e;
    ram_cell[    9753] = 32'h618d5c25;
    ram_cell[    9754] = 32'h3d5ca0f3;
    ram_cell[    9755] = 32'hce419acd;
    ram_cell[    9756] = 32'hc60d0ce1;
    ram_cell[    9757] = 32'h7c2cce42;
    ram_cell[    9758] = 32'h1973b336;
    ram_cell[    9759] = 32'h4111f6bc;
    ram_cell[    9760] = 32'ha11de84b;
    ram_cell[    9761] = 32'h0cfba25d;
    ram_cell[    9762] = 32'hee7565fb;
    ram_cell[    9763] = 32'hd5faeeef;
    ram_cell[    9764] = 32'h1d34050b;
    ram_cell[    9765] = 32'h43dd6596;
    ram_cell[    9766] = 32'h101acb47;
    ram_cell[    9767] = 32'ha033fadf;
    ram_cell[    9768] = 32'he99dba94;
    ram_cell[    9769] = 32'ha242d475;
    ram_cell[    9770] = 32'h891360c1;
    ram_cell[    9771] = 32'ha618a49a;
    ram_cell[    9772] = 32'ha278c2e7;
    ram_cell[    9773] = 32'h78da7364;
    ram_cell[    9774] = 32'ha455b70b;
    ram_cell[    9775] = 32'h9eea39f5;
    ram_cell[    9776] = 32'ha813f381;
    ram_cell[    9777] = 32'he22bcca2;
    ram_cell[    9778] = 32'hecd4ba3b;
    ram_cell[    9779] = 32'he10451dd;
    ram_cell[    9780] = 32'haf372720;
    ram_cell[    9781] = 32'h04ab667b;
    ram_cell[    9782] = 32'hfaf0aca7;
    ram_cell[    9783] = 32'h95767eb8;
    ram_cell[    9784] = 32'h58f8e410;
    ram_cell[    9785] = 32'h6826b0fa;
    ram_cell[    9786] = 32'h113bd74a;
    ram_cell[    9787] = 32'h88dcb130;
    ram_cell[    9788] = 32'ha561df32;
    ram_cell[    9789] = 32'h548e6540;
    ram_cell[    9790] = 32'h832771fb;
    ram_cell[    9791] = 32'h7084bcd9;
    ram_cell[    9792] = 32'h17f66e32;
    ram_cell[    9793] = 32'hb0ce8a1b;
    ram_cell[    9794] = 32'he025eb69;
    ram_cell[    9795] = 32'ha00282d9;
    ram_cell[    9796] = 32'h5491d268;
    ram_cell[    9797] = 32'hed00580c;
    ram_cell[    9798] = 32'heec621da;
    ram_cell[    9799] = 32'h23c59c0c;
    ram_cell[    9800] = 32'hdde0a7a8;
    ram_cell[    9801] = 32'h5de036ec;
    ram_cell[    9802] = 32'h78d4bacf;
    ram_cell[    9803] = 32'h67681810;
    ram_cell[    9804] = 32'hbae988d7;
    ram_cell[    9805] = 32'hf0272a8a;
    ram_cell[    9806] = 32'h8057c19e;
    ram_cell[    9807] = 32'hae420ae4;
    ram_cell[    9808] = 32'h9d408be1;
    ram_cell[    9809] = 32'heda82735;
    ram_cell[    9810] = 32'h89412293;
    ram_cell[    9811] = 32'hdca7dca3;
    ram_cell[    9812] = 32'h2b216484;
    ram_cell[    9813] = 32'hf753bf2c;
    ram_cell[    9814] = 32'h70800139;
    ram_cell[    9815] = 32'h9ecd9564;
    ram_cell[    9816] = 32'h215b17e8;
    ram_cell[    9817] = 32'h914d007c;
    ram_cell[    9818] = 32'h3843bbfa;
    ram_cell[    9819] = 32'h3e7fc012;
    ram_cell[    9820] = 32'heaad0f6d;
    ram_cell[    9821] = 32'h5bddcae9;
    ram_cell[    9822] = 32'he6797c66;
    ram_cell[    9823] = 32'h320fe3e0;
    ram_cell[    9824] = 32'hab14be8a;
    ram_cell[    9825] = 32'h66de2d54;
    ram_cell[    9826] = 32'he21c57f5;
    ram_cell[    9827] = 32'hc3aea141;
    ram_cell[    9828] = 32'h01dd775d;
    ram_cell[    9829] = 32'haf8bb1c0;
    ram_cell[    9830] = 32'h9ce2a260;
    ram_cell[    9831] = 32'h7be9b49e;
    ram_cell[    9832] = 32'hd50c1877;
    ram_cell[    9833] = 32'h73570092;
    ram_cell[    9834] = 32'h6c8dcad4;
    ram_cell[    9835] = 32'h960a7c24;
    ram_cell[    9836] = 32'h29d34675;
    ram_cell[    9837] = 32'hbd33c24d;
    ram_cell[    9838] = 32'h85489b9c;
    ram_cell[    9839] = 32'ha2d7ca48;
    ram_cell[    9840] = 32'h94ee62e8;
    ram_cell[    9841] = 32'h44177d1a;
    ram_cell[    9842] = 32'h730fa324;
    ram_cell[    9843] = 32'hd0c64016;
    ram_cell[    9844] = 32'h542b9e49;
    ram_cell[    9845] = 32'h228e04e1;
    ram_cell[    9846] = 32'hda445e67;
    ram_cell[    9847] = 32'h110f227f;
    ram_cell[    9848] = 32'h085b8568;
    ram_cell[    9849] = 32'h819eba09;
    ram_cell[    9850] = 32'h19c1d643;
    ram_cell[    9851] = 32'h8ed1c778;
    ram_cell[    9852] = 32'h9802c775;
    ram_cell[    9853] = 32'hc63fcc5c;
    ram_cell[    9854] = 32'h0773bd9b;
    ram_cell[    9855] = 32'h462cee5b;
    ram_cell[    9856] = 32'h77739987;
    ram_cell[    9857] = 32'h54231080;
    ram_cell[    9858] = 32'h95b3f6a3;
    ram_cell[    9859] = 32'h77c2a950;
    ram_cell[    9860] = 32'ha7dfd743;
    ram_cell[    9861] = 32'h5f3bbcff;
    ram_cell[    9862] = 32'h9efd9a48;
    ram_cell[    9863] = 32'hd7f4c0a6;
    ram_cell[    9864] = 32'h8149210e;
    ram_cell[    9865] = 32'h855347d2;
    ram_cell[    9866] = 32'h5e7cb0ae;
    ram_cell[    9867] = 32'h16d27249;
    ram_cell[    9868] = 32'h71e47b0f;
    ram_cell[    9869] = 32'hf4c9608f;
    ram_cell[    9870] = 32'h1ac97f56;
    ram_cell[    9871] = 32'ha682962a;
    ram_cell[    9872] = 32'he631bb7c;
    ram_cell[    9873] = 32'h501c46e1;
    ram_cell[    9874] = 32'hd1c8d193;
    ram_cell[    9875] = 32'h0543cd6e;
    ram_cell[    9876] = 32'h0b2a1c99;
    ram_cell[    9877] = 32'h9981d124;
    ram_cell[    9878] = 32'hbe0e0720;
    ram_cell[    9879] = 32'h14bcea41;
    ram_cell[    9880] = 32'hb7ae04eb;
    ram_cell[    9881] = 32'hd3fe7550;
    ram_cell[    9882] = 32'h62c56186;
    ram_cell[    9883] = 32'h492660d2;
    ram_cell[    9884] = 32'h2450c23e;
    ram_cell[    9885] = 32'hdb34d7da;
    ram_cell[    9886] = 32'hd9a074b7;
    ram_cell[    9887] = 32'hc421466a;
    ram_cell[    9888] = 32'h5e5d0919;
    ram_cell[    9889] = 32'h0e4aa30b;
    ram_cell[    9890] = 32'hf8e84ea4;
    ram_cell[    9891] = 32'h6938e6c3;
    ram_cell[    9892] = 32'h8f5e1a42;
    ram_cell[    9893] = 32'h6825dab3;
    ram_cell[    9894] = 32'hf19eb9e3;
    ram_cell[    9895] = 32'hf88964a5;
    ram_cell[    9896] = 32'h3a90f08d;
    ram_cell[    9897] = 32'hbb04a907;
    ram_cell[    9898] = 32'h5664c158;
    ram_cell[    9899] = 32'h4702b33c;
    ram_cell[    9900] = 32'h00502ae0;
    ram_cell[    9901] = 32'h967da105;
    ram_cell[    9902] = 32'h5f4df56f;
    ram_cell[    9903] = 32'h9c7e267b;
    ram_cell[    9904] = 32'h6adac23d;
    ram_cell[    9905] = 32'hda2b1b65;
    ram_cell[    9906] = 32'h6f2f6ec1;
    ram_cell[    9907] = 32'h91b30658;
    ram_cell[    9908] = 32'ha17fff85;
    ram_cell[    9909] = 32'ha11805cc;
    ram_cell[    9910] = 32'h7e79624a;
    ram_cell[    9911] = 32'hd6c67581;
    ram_cell[    9912] = 32'h395b69ed;
    ram_cell[    9913] = 32'h0fa14b9f;
    ram_cell[    9914] = 32'ha3ca8e8d;
    ram_cell[    9915] = 32'h49c94c9c;
    ram_cell[    9916] = 32'h0ade89b3;
    ram_cell[    9917] = 32'h2a286744;
    ram_cell[    9918] = 32'h9aff1485;
    ram_cell[    9919] = 32'h01e4f427;
    ram_cell[    9920] = 32'h8342cd6a;
    ram_cell[    9921] = 32'h72196e0d;
    ram_cell[    9922] = 32'h7fa65da0;
    ram_cell[    9923] = 32'h9a07e612;
    ram_cell[    9924] = 32'hec3ce6e1;
    ram_cell[    9925] = 32'h97e810be;
    ram_cell[    9926] = 32'h887287bf;
    ram_cell[    9927] = 32'h904347a0;
    ram_cell[    9928] = 32'h5641fa72;
    ram_cell[    9929] = 32'hf1b69edc;
    ram_cell[    9930] = 32'hf19e2498;
    ram_cell[    9931] = 32'h313a909b;
    ram_cell[    9932] = 32'h64263567;
    ram_cell[    9933] = 32'h4c477f0e;
    ram_cell[    9934] = 32'ha8e4319d;
    ram_cell[    9935] = 32'h31b61a0d;
    ram_cell[    9936] = 32'h84e59680;
    ram_cell[    9937] = 32'hb51521da;
    ram_cell[    9938] = 32'hc8a0ec35;
    ram_cell[    9939] = 32'h5fbccfd5;
    ram_cell[    9940] = 32'ha60893ed;
    ram_cell[    9941] = 32'ha243a28f;
    ram_cell[    9942] = 32'h8705bf64;
    ram_cell[    9943] = 32'h43c76843;
    ram_cell[    9944] = 32'h3b80c973;
    ram_cell[    9945] = 32'hc22a40e2;
    ram_cell[    9946] = 32'h5d3f9555;
    ram_cell[    9947] = 32'h5f343472;
    ram_cell[    9948] = 32'h639e5e38;
    ram_cell[    9949] = 32'hcdff7569;
    ram_cell[    9950] = 32'h818acb66;
    ram_cell[    9951] = 32'h82b94d4d;
    ram_cell[    9952] = 32'hd7f82eab;
    ram_cell[    9953] = 32'h6441660d;
    ram_cell[    9954] = 32'h426c0c78;
    ram_cell[    9955] = 32'h3ed02ee1;
    ram_cell[    9956] = 32'h339237fa;
    ram_cell[    9957] = 32'hedeaf08d;
    ram_cell[    9958] = 32'hfe68b5f9;
    ram_cell[    9959] = 32'h25ef8f84;
    ram_cell[    9960] = 32'hdccd39df;
    ram_cell[    9961] = 32'h588ddcbc;
    ram_cell[    9962] = 32'h4ac2c99c;
    ram_cell[    9963] = 32'h97603d43;
    ram_cell[    9964] = 32'hac131fbf;
    ram_cell[    9965] = 32'hb91e6ffa;
    ram_cell[    9966] = 32'he971a968;
    ram_cell[    9967] = 32'h637d5fea;
    ram_cell[    9968] = 32'h738ea09f;
    ram_cell[    9969] = 32'h65617861;
    ram_cell[    9970] = 32'h2ff20e04;
    ram_cell[    9971] = 32'h8ebd0b23;
    ram_cell[    9972] = 32'heda037e8;
    ram_cell[    9973] = 32'he5a09bf6;
    ram_cell[    9974] = 32'h17b39f03;
    ram_cell[    9975] = 32'hfc1d07b8;
    ram_cell[    9976] = 32'h6fbc346f;
    ram_cell[    9977] = 32'hff787ff4;
    ram_cell[    9978] = 32'hf2fde69f;
    ram_cell[    9979] = 32'hb532275c;
    ram_cell[    9980] = 32'hb01f5d83;
    ram_cell[    9981] = 32'h6e494259;
    ram_cell[    9982] = 32'h3c3fa32d;
    ram_cell[    9983] = 32'he5c44305;
    ram_cell[    9984] = 32'h7110cd70;
    ram_cell[    9985] = 32'h4f59c012;
    ram_cell[    9986] = 32'h8df416a4;
    ram_cell[    9987] = 32'hfa8cb536;
    ram_cell[    9988] = 32'hfe98db2a;
    ram_cell[    9989] = 32'h1030bc1c;
    ram_cell[    9990] = 32'hbd4e7086;
    ram_cell[    9991] = 32'h0313109e;
    ram_cell[    9992] = 32'h72ef7646;
    ram_cell[    9993] = 32'h53ad618b;
    ram_cell[    9994] = 32'h5ea2dc3f;
    ram_cell[    9995] = 32'h17c3d7b8;
    ram_cell[    9996] = 32'h0707f486;
    ram_cell[    9997] = 32'hbbb68a6d;
    ram_cell[    9998] = 32'h2267c242;
    ram_cell[    9999] = 32'h33fad173;
    ram_cell[   10000] = 32'h15e07ad6;
    ram_cell[   10001] = 32'he925f280;
    ram_cell[   10002] = 32'h3fc12887;
    ram_cell[   10003] = 32'hc2462e2c;
    ram_cell[   10004] = 32'h612af1c1;
    ram_cell[   10005] = 32'h390b6434;
    ram_cell[   10006] = 32'h05fe04ee;
    ram_cell[   10007] = 32'h6496c94e;
    ram_cell[   10008] = 32'hdb8e86ca;
    ram_cell[   10009] = 32'h69346ccc;
    ram_cell[   10010] = 32'h0bc90bf6;
    ram_cell[   10011] = 32'hb3098622;
    ram_cell[   10012] = 32'hd2366caa;
    ram_cell[   10013] = 32'h0a54bb3a;
    ram_cell[   10014] = 32'h2e5ddf05;
    ram_cell[   10015] = 32'hd29e1ce6;
    ram_cell[   10016] = 32'h22a05dba;
    ram_cell[   10017] = 32'h57f2b60a;
    ram_cell[   10018] = 32'h03931de4;
    ram_cell[   10019] = 32'hfba9791d;
    ram_cell[   10020] = 32'hc3cdf97b;
    ram_cell[   10021] = 32'h49498f10;
    ram_cell[   10022] = 32'h3799d75e;
    ram_cell[   10023] = 32'h7800beff;
    ram_cell[   10024] = 32'h33aae230;
    ram_cell[   10025] = 32'h0269dd14;
    ram_cell[   10026] = 32'h8877039c;
    ram_cell[   10027] = 32'h51025b4f;
    ram_cell[   10028] = 32'hb776bcf4;
    ram_cell[   10029] = 32'h09a272ca;
    ram_cell[   10030] = 32'h7d5b5485;
    ram_cell[   10031] = 32'h31d72f5d;
    ram_cell[   10032] = 32'he93316b4;
    ram_cell[   10033] = 32'h4e665abd;
    ram_cell[   10034] = 32'h78824b8f;
    ram_cell[   10035] = 32'h9927492b;
    ram_cell[   10036] = 32'h5d0bcb6b;
    ram_cell[   10037] = 32'ha62d56b4;
    ram_cell[   10038] = 32'h98e1facf;
    ram_cell[   10039] = 32'h8caaff94;
    ram_cell[   10040] = 32'ha1c0e243;
    ram_cell[   10041] = 32'h344ad1a3;
    ram_cell[   10042] = 32'h729883e7;
    ram_cell[   10043] = 32'he5407044;
    ram_cell[   10044] = 32'h2451500d;
    ram_cell[   10045] = 32'ha0ec524f;
    ram_cell[   10046] = 32'hef7d93f7;
    ram_cell[   10047] = 32'hdf68cf8e;
    ram_cell[   10048] = 32'h1545975b;
    ram_cell[   10049] = 32'h142f6292;
    ram_cell[   10050] = 32'h208e5c30;
    ram_cell[   10051] = 32'hb9fa138e;
    ram_cell[   10052] = 32'h70c3955b;
    ram_cell[   10053] = 32'h4db2a089;
    ram_cell[   10054] = 32'h60029c69;
    ram_cell[   10055] = 32'h32b5bc48;
    ram_cell[   10056] = 32'ha1fa969a;
    ram_cell[   10057] = 32'h1c51d89b;
    ram_cell[   10058] = 32'h2ec3ef83;
    ram_cell[   10059] = 32'hc2cc2d4d;
    ram_cell[   10060] = 32'h01acb066;
    ram_cell[   10061] = 32'h1636d44f;
    ram_cell[   10062] = 32'h0fc8b9ae;
    ram_cell[   10063] = 32'h21a7f37e;
    ram_cell[   10064] = 32'h4ea2a295;
    ram_cell[   10065] = 32'h1cad48a6;
    ram_cell[   10066] = 32'h3a87eb72;
    ram_cell[   10067] = 32'h91f77fe4;
    ram_cell[   10068] = 32'h197e62f6;
    ram_cell[   10069] = 32'he602027c;
    ram_cell[   10070] = 32'hb7911ccc;
    ram_cell[   10071] = 32'hff508634;
    ram_cell[   10072] = 32'h975511eb;
    ram_cell[   10073] = 32'haa0d19e3;
    ram_cell[   10074] = 32'hb65254c3;
    ram_cell[   10075] = 32'h31b8cf4c;
    ram_cell[   10076] = 32'h38266dd5;
    ram_cell[   10077] = 32'hfb04cb6d;
    ram_cell[   10078] = 32'h823397e1;
    ram_cell[   10079] = 32'hf94fe480;
    ram_cell[   10080] = 32'hc1dd6970;
    ram_cell[   10081] = 32'h1670eeab;
    ram_cell[   10082] = 32'hc94b5ff9;
    ram_cell[   10083] = 32'h99e06331;
    ram_cell[   10084] = 32'ha8dcc35c;
    ram_cell[   10085] = 32'hc16f06b7;
    ram_cell[   10086] = 32'h738211e3;
    ram_cell[   10087] = 32'hae62c844;
    ram_cell[   10088] = 32'h54f07b5f;
    ram_cell[   10089] = 32'he24f6b7b;
    ram_cell[   10090] = 32'h72c9e6df;
    ram_cell[   10091] = 32'h8162ce4b;
    ram_cell[   10092] = 32'h80435bb5;
    ram_cell[   10093] = 32'hd13a5e99;
    ram_cell[   10094] = 32'ha9103534;
    ram_cell[   10095] = 32'hc998d28f;
    ram_cell[   10096] = 32'h6b55f981;
    ram_cell[   10097] = 32'h9626cdd6;
    ram_cell[   10098] = 32'h8756e5ad;
    ram_cell[   10099] = 32'hecbed418;
    ram_cell[   10100] = 32'h96edadf8;
    ram_cell[   10101] = 32'h5eeaea1f;
    ram_cell[   10102] = 32'ha393a8c3;
    ram_cell[   10103] = 32'h15babbb6;
    ram_cell[   10104] = 32'h3ab2eee7;
    ram_cell[   10105] = 32'h54846dc1;
    ram_cell[   10106] = 32'h59f8015a;
    ram_cell[   10107] = 32'he628ebda;
    ram_cell[   10108] = 32'hdad7aed3;
    ram_cell[   10109] = 32'hd165ec01;
    ram_cell[   10110] = 32'hb78f5b31;
    ram_cell[   10111] = 32'hd3616116;
    ram_cell[   10112] = 32'h9ba34410;
    ram_cell[   10113] = 32'h4910477f;
    ram_cell[   10114] = 32'h71cb8cee;
    ram_cell[   10115] = 32'h598766f5;
    ram_cell[   10116] = 32'h0a1bb619;
    ram_cell[   10117] = 32'hb7d4ab5e;
    ram_cell[   10118] = 32'h36f6ae8b;
    ram_cell[   10119] = 32'h73a618ef;
    ram_cell[   10120] = 32'h4ed486a8;
    ram_cell[   10121] = 32'h4aca04f1;
    ram_cell[   10122] = 32'haa00f5af;
    ram_cell[   10123] = 32'hae072496;
    ram_cell[   10124] = 32'h7d6bba1f;
    ram_cell[   10125] = 32'h9ecbc767;
    ram_cell[   10126] = 32'h90490803;
    ram_cell[   10127] = 32'ha3770b84;
    ram_cell[   10128] = 32'h317755c8;
    ram_cell[   10129] = 32'hd1f5fa76;
    ram_cell[   10130] = 32'hdd0f6877;
    ram_cell[   10131] = 32'h5a2b46ad;
    ram_cell[   10132] = 32'h87c84c63;
    ram_cell[   10133] = 32'h4cc3f7c8;
    ram_cell[   10134] = 32'h520d2606;
    ram_cell[   10135] = 32'h3834ec8f;
    ram_cell[   10136] = 32'h0c4b8e79;
    ram_cell[   10137] = 32'h192288c1;
    ram_cell[   10138] = 32'h7d4f7423;
    ram_cell[   10139] = 32'h63905db4;
    ram_cell[   10140] = 32'hf8206e13;
    ram_cell[   10141] = 32'h542b9318;
    ram_cell[   10142] = 32'h2bf6565e;
    ram_cell[   10143] = 32'h5deebcac;
    ram_cell[   10144] = 32'hf81011db;
    ram_cell[   10145] = 32'h30ca8a28;
    ram_cell[   10146] = 32'hd4ecd2b4;
    ram_cell[   10147] = 32'h97265e09;
    ram_cell[   10148] = 32'hf1ed978c;
    ram_cell[   10149] = 32'h4d3beec1;
    ram_cell[   10150] = 32'h27691f4e;
    ram_cell[   10151] = 32'h5f556362;
    ram_cell[   10152] = 32'hca4881eb;
    ram_cell[   10153] = 32'h33c8d7e8;
    ram_cell[   10154] = 32'hbb1bae78;
    ram_cell[   10155] = 32'h63b07bd2;
    ram_cell[   10156] = 32'h6067fce1;
    ram_cell[   10157] = 32'h67588a51;
    ram_cell[   10158] = 32'hf7e74148;
    ram_cell[   10159] = 32'h8c708230;
    ram_cell[   10160] = 32'hdf623524;
    ram_cell[   10161] = 32'hf845a65e;
    ram_cell[   10162] = 32'h70994ee9;
    ram_cell[   10163] = 32'h39d92ce7;
    ram_cell[   10164] = 32'hed5d9bc3;
    ram_cell[   10165] = 32'hde5072e3;
    ram_cell[   10166] = 32'h33c5314e;
    ram_cell[   10167] = 32'h5664b035;
    ram_cell[   10168] = 32'hdea1da30;
    ram_cell[   10169] = 32'hb4645b08;
    ram_cell[   10170] = 32'hcb88be82;
    ram_cell[   10171] = 32'h0ca0df6b;
    ram_cell[   10172] = 32'h0f7be864;
    ram_cell[   10173] = 32'h631025b6;
    ram_cell[   10174] = 32'he6142662;
    ram_cell[   10175] = 32'hda2037f0;
    ram_cell[   10176] = 32'h37253d64;
    ram_cell[   10177] = 32'hb59f7dd7;
    ram_cell[   10178] = 32'h5998574a;
    ram_cell[   10179] = 32'hb3095d77;
    ram_cell[   10180] = 32'h7bde196a;
    ram_cell[   10181] = 32'hc79ca68a;
    ram_cell[   10182] = 32'ha1d1f05b;
    ram_cell[   10183] = 32'h3b82ed32;
    ram_cell[   10184] = 32'h3b8d2585;
    ram_cell[   10185] = 32'ha463d81d;
    ram_cell[   10186] = 32'h2fb9b24f;
    ram_cell[   10187] = 32'h730785fc;
    ram_cell[   10188] = 32'hddc69e4a;
    ram_cell[   10189] = 32'hf540102d;
    ram_cell[   10190] = 32'h6f90cd85;
    ram_cell[   10191] = 32'h9171a217;
    ram_cell[   10192] = 32'h967fac6b;
    ram_cell[   10193] = 32'hc89d0b23;
    ram_cell[   10194] = 32'h85dde18e;
    ram_cell[   10195] = 32'h35fc8c72;
    ram_cell[   10196] = 32'h4ae43d2a;
    ram_cell[   10197] = 32'h204ff6ee;
    ram_cell[   10198] = 32'h084c0afc;
    ram_cell[   10199] = 32'hd12bb314;
    ram_cell[   10200] = 32'h4fdde625;
    ram_cell[   10201] = 32'h8bd7dacb;
    ram_cell[   10202] = 32'h6122242b;
    ram_cell[   10203] = 32'hd537f869;
    ram_cell[   10204] = 32'h57485edb;
    ram_cell[   10205] = 32'h70bda6d0;
    ram_cell[   10206] = 32'h9903a6e2;
    ram_cell[   10207] = 32'hf90f0e93;
    ram_cell[   10208] = 32'he603e855;
    ram_cell[   10209] = 32'h3647a1f6;
    ram_cell[   10210] = 32'hc9de528e;
    ram_cell[   10211] = 32'h34309f68;
    ram_cell[   10212] = 32'h5a9a1d0c;
    ram_cell[   10213] = 32'h01423dbf;
    ram_cell[   10214] = 32'h9f78d54f;
    ram_cell[   10215] = 32'hb00e7621;
    ram_cell[   10216] = 32'hd67d00b1;
    ram_cell[   10217] = 32'h86d43d38;
    ram_cell[   10218] = 32'h12352c22;
    ram_cell[   10219] = 32'he62ea442;
    ram_cell[   10220] = 32'h04240e9b;
    ram_cell[   10221] = 32'hef0a796a;
    ram_cell[   10222] = 32'hcbaa2d8e;
    ram_cell[   10223] = 32'hc0a312b4;
    ram_cell[   10224] = 32'h44decd42;
    ram_cell[   10225] = 32'hb1736e5a;
    ram_cell[   10226] = 32'h1cc41ddc;
    ram_cell[   10227] = 32'hcc35f18d;
    ram_cell[   10228] = 32'h11379f3f;
    ram_cell[   10229] = 32'hf29b0295;
    ram_cell[   10230] = 32'h119d1041;
    ram_cell[   10231] = 32'h432c2921;
    ram_cell[   10232] = 32'h7637b78e;
    ram_cell[   10233] = 32'hcadae4c3;
    ram_cell[   10234] = 32'h9d28d702;
    ram_cell[   10235] = 32'h0b19bc07;
    ram_cell[   10236] = 32'h7ba96484;
    ram_cell[   10237] = 32'h96c07f03;
    ram_cell[   10238] = 32'h35653bc8;
    ram_cell[   10239] = 32'h9fa9b021;
    ram_cell[   10240] = 32'hf00669c5;
    ram_cell[   10241] = 32'h9e0cfb7d;
    ram_cell[   10242] = 32'hb18ea4a0;
    ram_cell[   10243] = 32'h789d7898;
    ram_cell[   10244] = 32'h01585e82;
    ram_cell[   10245] = 32'h307b6aa8;
    ram_cell[   10246] = 32'h29482030;
    ram_cell[   10247] = 32'h7687c163;
    ram_cell[   10248] = 32'h28c6a111;
    ram_cell[   10249] = 32'hfda78b00;
    ram_cell[   10250] = 32'hf4c2497e;
    ram_cell[   10251] = 32'h5fb712ce;
    ram_cell[   10252] = 32'h5a77cdde;
    ram_cell[   10253] = 32'h7c5627d8;
    ram_cell[   10254] = 32'h69b0b6c1;
    ram_cell[   10255] = 32'h1f15cd41;
    ram_cell[   10256] = 32'hdacd6097;
    ram_cell[   10257] = 32'ha7c50f03;
    ram_cell[   10258] = 32'h20885c64;
    ram_cell[   10259] = 32'h28778fef;
    ram_cell[   10260] = 32'h1cf744e2;
    ram_cell[   10261] = 32'h2ac8e06d;
    ram_cell[   10262] = 32'h3ac33c0d;
    ram_cell[   10263] = 32'h03c1967e;
    ram_cell[   10264] = 32'heac577a8;
    ram_cell[   10265] = 32'hc8a4af3f;
    ram_cell[   10266] = 32'h5218dffa;
    ram_cell[   10267] = 32'had23c21b;
    ram_cell[   10268] = 32'h68ba397b;
    ram_cell[   10269] = 32'h29de54ca;
    ram_cell[   10270] = 32'h4cda5ffe;
    ram_cell[   10271] = 32'hd4631f50;
    ram_cell[   10272] = 32'h07f53e51;
    ram_cell[   10273] = 32'h2b7549a3;
    ram_cell[   10274] = 32'h144dd729;
    ram_cell[   10275] = 32'hf9709d2e;
    ram_cell[   10276] = 32'h10e76f45;
    ram_cell[   10277] = 32'had04102c;
    ram_cell[   10278] = 32'hf4b37491;
    ram_cell[   10279] = 32'h25c94a4e;
    ram_cell[   10280] = 32'hd0477019;
    ram_cell[   10281] = 32'hf16e2c21;
    ram_cell[   10282] = 32'h7efc2701;
    ram_cell[   10283] = 32'hf3139f14;
    ram_cell[   10284] = 32'hca09266f;
    ram_cell[   10285] = 32'h305c472b;
    ram_cell[   10286] = 32'hee37d436;
    ram_cell[   10287] = 32'hcc7c36d4;
    ram_cell[   10288] = 32'h4078a4d4;
    ram_cell[   10289] = 32'h4616609d;
    ram_cell[   10290] = 32'h0cb31171;
    ram_cell[   10291] = 32'h9005d7e8;
    ram_cell[   10292] = 32'hac83d1f9;
    ram_cell[   10293] = 32'h756c1a43;
    ram_cell[   10294] = 32'h8f9e63bb;
    ram_cell[   10295] = 32'heab85d3d;
    ram_cell[   10296] = 32'h6f10916a;
    ram_cell[   10297] = 32'h0abb4053;
    ram_cell[   10298] = 32'h74a592fc;
    ram_cell[   10299] = 32'h3bb3bb5f;
    ram_cell[   10300] = 32'h7b32275c;
    ram_cell[   10301] = 32'h20e1fc91;
    ram_cell[   10302] = 32'h055989d8;
    ram_cell[   10303] = 32'he51d4584;
    ram_cell[   10304] = 32'h68f1db93;
    ram_cell[   10305] = 32'hc5dd4d7f;
    ram_cell[   10306] = 32'h3f59f139;
    ram_cell[   10307] = 32'h5348360f;
    ram_cell[   10308] = 32'hbe95e840;
    ram_cell[   10309] = 32'h76e73a69;
    ram_cell[   10310] = 32'h4742af6a;
    ram_cell[   10311] = 32'h71d4ddab;
    ram_cell[   10312] = 32'hab8c3677;
    ram_cell[   10313] = 32'h35b21a71;
    ram_cell[   10314] = 32'hec764a8f;
    ram_cell[   10315] = 32'h690a60d7;
    ram_cell[   10316] = 32'h1317cc52;
    ram_cell[   10317] = 32'he035e758;
    ram_cell[   10318] = 32'hcb45c1bf;
    ram_cell[   10319] = 32'h25dc2576;
    ram_cell[   10320] = 32'h44cc78eb;
    ram_cell[   10321] = 32'h757c5c06;
    ram_cell[   10322] = 32'h2a5f7ebe;
    ram_cell[   10323] = 32'h74e50296;
    ram_cell[   10324] = 32'h179517d5;
    ram_cell[   10325] = 32'h8f7685f9;
    ram_cell[   10326] = 32'hfaed2aa3;
    ram_cell[   10327] = 32'h1aaf50f1;
    ram_cell[   10328] = 32'hd216fc6c;
    ram_cell[   10329] = 32'h44ec7876;
    ram_cell[   10330] = 32'h1a9fb901;
    ram_cell[   10331] = 32'h64fedfb9;
    ram_cell[   10332] = 32'h00a5e66d;
    ram_cell[   10333] = 32'h2cca2969;
    ram_cell[   10334] = 32'h75834883;
    ram_cell[   10335] = 32'hb819dc45;
    ram_cell[   10336] = 32'hb832d177;
    ram_cell[   10337] = 32'h53514f0a;
    ram_cell[   10338] = 32'ha737bb36;
    ram_cell[   10339] = 32'h05898ba9;
    ram_cell[   10340] = 32'h0d38b287;
    ram_cell[   10341] = 32'hdf9d4333;
    ram_cell[   10342] = 32'hfb4280a9;
    ram_cell[   10343] = 32'h6661482a;
    ram_cell[   10344] = 32'hb3a64a20;
    ram_cell[   10345] = 32'h48eef46e;
    ram_cell[   10346] = 32'hd30871b6;
    ram_cell[   10347] = 32'h8b819376;
    ram_cell[   10348] = 32'h71457477;
    ram_cell[   10349] = 32'h063c38bc;
    ram_cell[   10350] = 32'hfbcee2c8;
    ram_cell[   10351] = 32'h13611c84;
    ram_cell[   10352] = 32'h260a0d49;
    ram_cell[   10353] = 32'h7a2769a2;
    ram_cell[   10354] = 32'h3b7d1be2;
    ram_cell[   10355] = 32'haeff59e5;
    ram_cell[   10356] = 32'hdf405228;
    ram_cell[   10357] = 32'h7b375767;
    ram_cell[   10358] = 32'h82094878;
    ram_cell[   10359] = 32'h4a66d909;
    ram_cell[   10360] = 32'h68957b5d;
    ram_cell[   10361] = 32'h87cfa84e;
    ram_cell[   10362] = 32'h23bde6a3;
    ram_cell[   10363] = 32'h6e28b0ee;
    ram_cell[   10364] = 32'h7311e145;
    ram_cell[   10365] = 32'h49aaab80;
    ram_cell[   10366] = 32'h6424b23c;
    ram_cell[   10367] = 32'hf8036181;
    ram_cell[   10368] = 32'h3b272e2b;
    ram_cell[   10369] = 32'hfa4fe138;
    ram_cell[   10370] = 32'hdf54a050;
    ram_cell[   10371] = 32'h117dbd7e;
    ram_cell[   10372] = 32'h4c7a1a75;
    ram_cell[   10373] = 32'h49a0f3d7;
    ram_cell[   10374] = 32'hd90fcd65;
    ram_cell[   10375] = 32'h9fb8b813;
    ram_cell[   10376] = 32'h852fa639;
    ram_cell[   10377] = 32'he526dbe0;
    ram_cell[   10378] = 32'h075848d5;
    ram_cell[   10379] = 32'h76d64a1c;
    ram_cell[   10380] = 32'h92d2ef6f;
    ram_cell[   10381] = 32'h1b38ccb3;
    ram_cell[   10382] = 32'h2b9d9148;
    ram_cell[   10383] = 32'h7c318214;
    ram_cell[   10384] = 32'h47305208;
    ram_cell[   10385] = 32'haffb7b58;
    ram_cell[   10386] = 32'h8cd809f9;
    ram_cell[   10387] = 32'hf799a46c;
    ram_cell[   10388] = 32'ha4bef92a;
    ram_cell[   10389] = 32'h0dbb40bb;
    ram_cell[   10390] = 32'h8166f83a;
    ram_cell[   10391] = 32'ha9ca8df5;
    ram_cell[   10392] = 32'h5ff519f6;
    ram_cell[   10393] = 32'h159722f7;
    ram_cell[   10394] = 32'h419a352d;
    ram_cell[   10395] = 32'hcafe656b;
    ram_cell[   10396] = 32'h92688051;
    ram_cell[   10397] = 32'hdbede5d7;
    ram_cell[   10398] = 32'hac1b7ecc;
    ram_cell[   10399] = 32'h2cc74fde;
    ram_cell[   10400] = 32'he9d75516;
    ram_cell[   10401] = 32'h8a006302;
    ram_cell[   10402] = 32'h836da2c0;
    ram_cell[   10403] = 32'h5d1d2e0b;
    ram_cell[   10404] = 32'he644deb0;
    ram_cell[   10405] = 32'hd00550eb;
    ram_cell[   10406] = 32'hba64a56b;
    ram_cell[   10407] = 32'h38dd3871;
    ram_cell[   10408] = 32'hcdb2bb22;
    ram_cell[   10409] = 32'h7951f663;
    ram_cell[   10410] = 32'heee4eebd;
    ram_cell[   10411] = 32'h81738960;
    ram_cell[   10412] = 32'h53972ae3;
    ram_cell[   10413] = 32'h116deeb1;
    ram_cell[   10414] = 32'h62184f15;
    ram_cell[   10415] = 32'h95e7012e;
    ram_cell[   10416] = 32'h7058e799;
    ram_cell[   10417] = 32'h390629b3;
    ram_cell[   10418] = 32'h998cd48b;
    ram_cell[   10419] = 32'h1a58dac6;
    ram_cell[   10420] = 32'h13aef940;
    ram_cell[   10421] = 32'hd6bc2c42;
    ram_cell[   10422] = 32'h94560417;
    ram_cell[   10423] = 32'h171f6205;
    ram_cell[   10424] = 32'h2a61ba3a;
    ram_cell[   10425] = 32'h05d88195;
    ram_cell[   10426] = 32'h75bc0ca3;
    ram_cell[   10427] = 32'h00d22167;
    ram_cell[   10428] = 32'h36f4da4e;
    ram_cell[   10429] = 32'h5d6ba450;
    ram_cell[   10430] = 32'hc87af082;
    ram_cell[   10431] = 32'ha11fda0e;
    ram_cell[   10432] = 32'h4aa000e3;
    ram_cell[   10433] = 32'h751d0418;
    ram_cell[   10434] = 32'hd6e46196;
    ram_cell[   10435] = 32'hb3a3905a;
    ram_cell[   10436] = 32'h67b6b0fa;
    ram_cell[   10437] = 32'h77717833;
    ram_cell[   10438] = 32'h9481a4f3;
    ram_cell[   10439] = 32'hf0c84f59;
    ram_cell[   10440] = 32'h6328bffd;
    ram_cell[   10441] = 32'hbceaf70e;
    ram_cell[   10442] = 32'hb0d5392b;
    ram_cell[   10443] = 32'h2eb0a871;
    ram_cell[   10444] = 32'h14593f77;
    ram_cell[   10445] = 32'h9ccc134c;
    ram_cell[   10446] = 32'h8288339d;
    ram_cell[   10447] = 32'h43fe5fb9;
    ram_cell[   10448] = 32'h9a465f01;
    ram_cell[   10449] = 32'h2cf8b0f8;
    ram_cell[   10450] = 32'h150c0cea;
    ram_cell[   10451] = 32'hd938b027;
    ram_cell[   10452] = 32'h66c3ed0b;
    ram_cell[   10453] = 32'he58ab2f9;
    ram_cell[   10454] = 32'h7a3c3390;
    ram_cell[   10455] = 32'h1fb8611f;
    ram_cell[   10456] = 32'hb1046dd0;
    ram_cell[   10457] = 32'hdd36ada5;
    ram_cell[   10458] = 32'h6042418c;
    ram_cell[   10459] = 32'h80b2fa80;
    ram_cell[   10460] = 32'h1ddf619b;
    ram_cell[   10461] = 32'h54853d98;
    ram_cell[   10462] = 32'he7967f12;
    ram_cell[   10463] = 32'hd97e6112;
    ram_cell[   10464] = 32'h0a819c65;
    ram_cell[   10465] = 32'hf7891402;
    ram_cell[   10466] = 32'h4889f178;
    ram_cell[   10467] = 32'h7d59e530;
    ram_cell[   10468] = 32'heffea037;
    ram_cell[   10469] = 32'h1a0701b7;
    ram_cell[   10470] = 32'h0621bbb1;
    ram_cell[   10471] = 32'hfb122e14;
    ram_cell[   10472] = 32'h8ec7bf7d;
    ram_cell[   10473] = 32'h93c22b0d;
    ram_cell[   10474] = 32'h92bef918;
    ram_cell[   10475] = 32'hc2f2be03;
    ram_cell[   10476] = 32'h9ec8e768;
    ram_cell[   10477] = 32'h2669d4b5;
    ram_cell[   10478] = 32'h4055190b;
    ram_cell[   10479] = 32'h093cc5d3;
    ram_cell[   10480] = 32'h320a0875;
    ram_cell[   10481] = 32'ha3150ae4;
    ram_cell[   10482] = 32'h217b6dee;
    ram_cell[   10483] = 32'hdd7ca5d3;
    ram_cell[   10484] = 32'h7085014f;
    ram_cell[   10485] = 32'h44fb463c;
    ram_cell[   10486] = 32'hb9f361db;
    ram_cell[   10487] = 32'h2a0b5409;
    ram_cell[   10488] = 32'hed6a329b;
    ram_cell[   10489] = 32'he64fc6cf;
    ram_cell[   10490] = 32'h80554437;
    ram_cell[   10491] = 32'h34ce1531;
    ram_cell[   10492] = 32'h98f4b3b9;
    ram_cell[   10493] = 32'h2a86fd9d;
    ram_cell[   10494] = 32'ha90743bf;
    ram_cell[   10495] = 32'hcce59b8d;
    ram_cell[   10496] = 32'h98c97f53;
    ram_cell[   10497] = 32'h80fb96de;
    ram_cell[   10498] = 32'hda9b734d;
    ram_cell[   10499] = 32'h3b2ba358;
    ram_cell[   10500] = 32'hc75f30bb;
    ram_cell[   10501] = 32'hf463d385;
    ram_cell[   10502] = 32'heb5311c9;
    ram_cell[   10503] = 32'h9842693e;
    ram_cell[   10504] = 32'hdb71c42d;
    ram_cell[   10505] = 32'h53b4972d;
    ram_cell[   10506] = 32'h393d6a0d;
    ram_cell[   10507] = 32'h80bba72c;
    ram_cell[   10508] = 32'hbf756f1d;
    ram_cell[   10509] = 32'h1a6b220d;
    ram_cell[   10510] = 32'h4511f0a0;
    ram_cell[   10511] = 32'h38d39655;
    ram_cell[   10512] = 32'he4a2d7ed;
    ram_cell[   10513] = 32'h910a317f;
    ram_cell[   10514] = 32'h50d3702f;
    ram_cell[   10515] = 32'h1ec9035c;
    ram_cell[   10516] = 32'h49dc0aaf;
    ram_cell[   10517] = 32'he29c4449;
    ram_cell[   10518] = 32'h26e93327;
    ram_cell[   10519] = 32'h47d80b57;
    ram_cell[   10520] = 32'h8fc67f5b;
    ram_cell[   10521] = 32'h8c7221dc;
    ram_cell[   10522] = 32'hbfdbb696;
    ram_cell[   10523] = 32'h037b7ab1;
    ram_cell[   10524] = 32'h4958f586;
    ram_cell[   10525] = 32'h78330140;
    ram_cell[   10526] = 32'h7b58ceba;
    ram_cell[   10527] = 32'h4bf389c3;
    ram_cell[   10528] = 32'h93102722;
    ram_cell[   10529] = 32'hd840c1fc;
    ram_cell[   10530] = 32'h6a301c03;
    ram_cell[   10531] = 32'h290022aa;
    ram_cell[   10532] = 32'h1324b4de;
    ram_cell[   10533] = 32'hc3cb2348;
    ram_cell[   10534] = 32'ha238f4f7;
    ram_cell[   10535] = 32'h990dc6e9;
    ram_cell[   10536] = 32'hf32b3ca6;
    ram_cell[   10537] = 32'h49e9a44d;
    ram_cell[   10538] = 32'hb4af5707;
    ram_cell[   10539] = 32'hd307d19e;
    ram_cell[   10540] = 32'h74d90ad6;
    ram_cell[   10541] = 32'h1a1c58b4;
    ram_cell[   10542] = 32'ha442c637;
    ram_cell[   10543] = 32'h74291a7c;
    ram_cell[   10544] = 32'h64e110f2;
    ram_cell[   10545] = 32'h6972786e;
    ram_cell[   10546] = 32'h6d5f1202;
    ram_cell[   10547] = 32'h816a1bfd;
    ram_cell[   10548] = 32'hec4b6919;
    ram_cell[   10549] = 32'hffd845ef;
    ram_cell[   10550] = 32'h983462c6;
    ram_cell[   10551] = 32'he4f24c2e;
    ram_cell[   10552] = 32'hfcb93dcb;
    ram_cell[   10553] = 32'h1679a3ce;
    ram_cell[   10554] = 32'hd35a9735;
    ram_cell[   10555] = 32'h7597a4b9;
    ram_cell[   10556] = 32'h35b901e8;
    ram_cell[   10557] = 32'h8bda9ee2;
    ram_cell[   10558] = 32'h7b2ac460;
    ram_cell[   10559] = 32'he4726463;
    ram_cell[   10560] = 32'h40518e2e;
    ram_cell[   10561] = 32'h9754a977;
    ram_cell[   10562] = 32'hc90bcedc;
    ram_cell[   10563] = 32'h4466a372;
    ram_cell[   10564] = 32'h352619dd;
    ram_cell[   10565] = 32'hfeb5865f;
    ram_cell[   10566] = 32'h5f9849fa;
    ram_cell[   10567] = 32'h713ea697;
    ram_cell[   10568] = 32'h045984ed;
    ram_cell[   10569] = 32'h53eb801e;
    ram_cell[   10570] = 32'h38afe676;
    ram_cell[   10571] = 32'h6beed24d;
    ram_cell[   10572] = 32'h15511a69;
    ram_cell[   10573] = 32'hd18a6b09;
    ram_cell[   10574] = 32'h00578b19;
    ram_cell[   10575] = 32'ha2f947da;
    ram_cell[   10576] = 32'h7a9e9f48;
    ram_cell[   10577] = 32'h72f7074c;
    ram_cell[   10578] = 32'h037b78d0;
    ram_cell[   10579] = 32'h74343936;
    ram_cell[   10580] = 32'h6f5617a3;
    ram_cell[   10581] = 32'ha1f34c19;
    ram_cell[   10582] = 32'h4f1e2094;
    ram_cell[   10583] = 32'h76c181d4;
    ram_cell[   10584] = 32'h00cc9e0d;
    ram_cell[   10585] = 32'h7f7f4745;
    ram_cell[   10586] = 32'h6bfe462d;
    ram_cell[   10587] = 32'hcd9bf5f9;
    ram_cell[   10588] = 32'hda93a638;
    ram_cell[   10589] = 32'h60c68fee;
    ram_cell[   10590] = 32'h11e33b25;
    ram_cell[   10591] = 32'h4e892e9d;
    ram_cell[   10592] = 32'h84149aca;
    ram_cell[   10593] = 32'hbe7443fd;
    ram_cell[   10594] = 32'h9d1b0ac2;
    ram_cell[   10595] = 32'h5c6f5c31;
    ram_cell[   10596] = 32'he26eff30;
    ram_cell[   10597] = 32'h0d363841;
    ram_cell[   10598] = 32'ha658acd4;
    ram_cell[   10599] = 32'h1b994b55;
    ram_cell[   10600] = 32'hccd2f5ba;
    ram_cell[   10601] = 32'h636fed80;
    ram_cell[   10602] = 32'h2e9100c4;
    ram_cell[   10603] = 32'h3d2305e6;
    ram_cell[   10604] = 32'hf6918f57;
    ram_cell[   10605] = 32'h16386a37;
    ram_cell[   10606] = 32'hc76d2917;
    ram_cell[   10607] = 32'hdca9ea5a;
    ram_cell[   10608] = 32'haa578273;
    ram_cell[   10609] = 32'h4f2d9da3;
    ram_cell[   10610] = 32'h2ecaa0ad;
    ram_cell[   10611] = 32'h8a06200a;
    ram_cell[   10612] = 32'h82bf1fbc;
    ram_cell[   10613] = 32'h7590a6b7;
    ram_cell[   10614] = 32'h35c4ffdb;
    ram_cell[   10615] = 32'h5332fdc6;
    ram_cell[   10616] = 32'h80d16ced;
    ram_cell[   10617] = 32'h7175dccd;
    ram_cell[   10618] = 32'h248e2480;
    ram_cell[   10619] = 32'h89fb77af;
    ram_cell[   10620] = 32'h1cbeaaa9;
    ram_cell[   10621] = 32'h1a28bf57;
    ram_cell[   10622] = 32'h81808917;
    ram_cell[   10623] = 32'h1a71d7b6;
    ram_cell[   10624] = 32'h6b8148d0;
    ram_cell[   10625] = 32'h14e40cba;
    ram_cell[   10626] = 32'h4bc52bb6;
    ram_cell[   10627] = 32'h369f97cc;
    ram_cell[   10628] = 32'h3d83bfd7;
    ram_cell[   10629] = 32'h003940b2;
    ram_cell[   10630] = 32'h9bd57bf8;
    ram_cell[   10631] = 32'h60fa31e4;
    ram_cell[   10632] = 32'ha9daf487;
    ram_cell[   10633] = 32'h2d71a7ce;
    ram_cell[   10634] = 32'he486bfa4;
    ram_cell[   10635] = 32'h1f081652;
    ram_cell[   10636] = 32'h9184575d;
    ram_cell[   10637] = 32'h9129c795;
    ram_cell[   10638] = 32'h9f7e5b7e;
    ram_cell[   10639] = 32'he6f53b72;
    ram_cell[   10640] = 32'hb8db426c;
    ram_cell[   10641] = 32'hffed7824;
    ram_cell[   10642] = 32'haa7da86a;
    ram_cell[   10643] = 32'h68949638;
    ram_cell[   10644] = 32'hed66bedf;
    ram_cell[   10645] = 32'h1e6adeb8;
    ram_cell[   10646] = 32'h219b0703;
    ram_cell[   10647] = 32'hb28f69c3;
    ram_cell[   10648] = 32'h8050c87a;
    ram_cell[   10649] = 32'hd4df55ef;
    ram_cell[   10650] = 32'h3c487f70;
    ram_cell[   10651] = 32'h700baea6;
    ram_cell[   10652] = 32'h415be583;
    ram_cell[   10653] = 32'h7712b4d1;
    ram_cell[   10654] = 32'h3234094e;
    ram_cell[   10655] = 32'hb4398ed5;
    ram_cell[   10656] = 32'h84dbad00;
    ram_cell[   10657] = 32'he13e8efd;
    ram_cell[   10658] = 32'h74af0bff;
    ram_cell[   10659] = 32'hbd01d9b3;
    ram_cell[   10660] = 32'h56656a2a;
    ram_cell[   10661] = 32'hc984fbf7;
    ram_cell[   10662] = 32'h456d35e8;
    ram_cell[   10663] = 32'h1856ed67;
    ram_cell[   10664] = 32'h38c32958;
    ram_cell[   10665] = 32'h3e2d5009;
    ram_cell[   10666] = 32'h8fd3ba38;
    ram_cell[   10667] = 32'ha49094fb;
    ram_cell[   10668] = 32'hd39b6907;
    ram_cell[   10669] = 32'h8196473d;
    ram_cell[   10670] = 32'hc213ec06;
    ram_cell[   10671] = 32'h5c46e08a;
    ram_cell[   10672] = 32'h23745f0b;
    ram_cell[   10673] = 32'h833e7d9f;
    ram_cell[   10674] = 32'hc2f25e76;
    ram_cell[   10675] = 32'h4c7ae1fa;
    ram_cell[   10676] = 32'h59fc39d5;
    ram_cell[   10677] = 32'h9e6745b1;
    ram_cell[   10678] = 32'headeb24e;
    ram_cell[   10679] = 32'h437226f7;
    ram_cell[   10680] = 32'h97d25de7;
    ram_cell[   10681] = 32'h0aac961d;
    ram_cell[   10682] = 32'h89bccb46;
    ram_cell[   10683] = 32'h1aedf562;
    ram_cell[   10684] = 32'h504e1abd;
    ram_cell[   10685] = 32'h103f4ec8;
    ram_cell[   10686] = 32'h6f1129ce;
    ram_cell[   10687] = 32'h91b4852c;
    ram_cell[   10688] = 32'h6b414530;
    ram_cell[   10689] = 32'h66089df6;
    ram_cell[   10690] = 32'h23251b94;
    ram_cell[   10691] = 32'h0fe99b3e;
    ram_cell[   10692] = 32'h25afe1b9;
    ram_cell[   10693] = 32'h02ab6c9f;
    ram_cell[   10694] = 32'h0d89e26b;
    ram_cell[   10695] = 32'hef146f45;
    ram_cell[   10696] = 32'hec90b36e;
    ram_cell[   10697] = 32'h91826216;
    ram_cell[   10698] = 32'h3b5d60a3;
    ram_cell[   10699] = 32'hfab0ac3d;
    ram_cell[   10700] = 32'ha75bbf31;
    ram_cell[   10701] = 32'h70403c22;
    ram_cell[   10702] = 32'had2b6387;
    ram_cell[   10703] = 32'h9ea44f10;
    ram_cell[   10704] = 32'h3b743cf8;
    ram_cell[   10705] = 32'h72f72a84;
    ram_cell[   10706] = 32'hbdad1c3f;
    ram_cell[   10707] = 32'hb3ac6578;
    ram_cell[   10708] = 32'h4e1ba7ea;
    ram_cell[   10709] = 32'h873a32d6;
    ram_cell[   10710] = 32'haa76589e;
    ram_cell[   10711] = 32'h79586587;
    ram_cell[   10712] = 32'hdafa01df;
    ram_cell[   10713] = 32'h4c63f264;
    ram_cell[   10714] = 32'he74873d6;
    ram_cell[   10715] = 32'h0311bf96;
    ram_cell[   10716] = 32'h958c75e5;
    ram_cell[   10717] = 32'h0a98cf24;
    ram_cell[   10718] = 32'h09a70dc3;
    ram_cell[   10719] = 32'h9f4ac419;
    ram_cell[   10720] = 32'h855cc736;
    ram_cell[   10721] = 32'h48a7501c;
    ram_cell[   10722] = 32'h58bfb3e2;
    ram_cell[   10723] = 32'he48d9da8;
    ram_cell[   10724] = 32'h8e119b4f;
    ram_cell[   10725] = 32'hb2b752de;
    ram_cell[   10726] = 32'h57dec7cd;
    ram_cell[   10727] = 32'hefd38495;
    ram_cell[   10728] = 32'h3475b798;
    ram_cell[   10729] = 32'h8dbcadd0;
    ram_cell[   10730] = 32'h523bef1b;
    ram_cell[   10731] = 32'h0f87c89c;
    ram_cell[   10732] = 32'h4333dcec;
    ram_cell[   10733] = 32'h1f95ce3d;
    ram_cell[   10734] = 32'h0f36a718;
    ram_cell[   10735] = 32'h329620a6;
    ram_cell[   10736] = 32'h9c221046;
    ram_cell[   10737] = 32'h936eeeea;
    ram_cell[   10738] = 32'h64fadd1b;
    ram_cell[   10739] = 32'hbae64a54;
    ram_cell[   10740] = 32'h6cc078ca;
    ram_cell[   10741] = 32'hf662797c;
    ram_cell[   10742] = 32'h4633a99e;
    ram_cell[   10743] = 32'h47a6489b;
    ram_cell[   10744] = 32'h7c51209a;
    ram_cell[   10745] = 32'h3954a825;
    ram_cell[   10746] = 32'hd24ff072;
    ram_cell[   10747] = 32'hc4e5fc4c;
    ram_cell[   10748] = 32'hf65618ed;
    ram_cell[   10749] = 32'h9288af2b;
    ram_cell[   10750] = 32'h645265e3;
    ram_cell[   10751] = 32'hb52ba882;
    ram_cell[   10752] = 32'h9e549e8c;
    ram_cell[   10753] = 32'hcb656000;
    ram_cell[   10754] = 32'h5ef1e3de;
    ram_cell[   10755] = 32'h8952c563;
    ram_cell[   10756] = 32'h9711d38c;
    ram_cell[   10757] = 32'h1e96b55a;
    ram_cell[   10758] = 32'hc62a2359;
    ram_cell[   10759] = 32'h4b59727f;
    ram_cell[   10760] = 32'hbd130db4;
    ram_cell[   10761] = 32'h62cfc3a7;
    ram_cell[   10762] = 32'h220cccc1;
    ram_cell[   10763] = 32'h4edb1bbb;
    ram_cell[   10764] = 32'hb7b8f519;
    ram_cell[   10765] = 32'h30c138f6;
    ram_cell[   10766] = 32'h6650f17b;
    ram_cell[   10767] = 32'hd728f91e;
    ram_cell[   10768] = 32'h76844afb;
    ram_cell[   10769] = 32'h3924fa9b;
    ram_cell[   10770] = 32'h076b5c82;
    ram_cell[   10771] = 32'hb39b185c;
    ram_cell[   10772] = 32'ha84aa605;
    ram_cell[   10773] = 32'hf5556bc3;
    ram_cell[   10774] = 32'h80a25829;
    ram_cell[   10775] = 32'hb9d102d7;
    ram_cell[   10776] = 32'h2e771933;
    ram_cell[   10777] = 32'h30440df0;
    ram_cell[   10778] = 32'hb7cabf20;
    ram_cell[   10779] = 32'h9522769f;
    ram_cell[   10780] = 32'hcd474577;
    ram_cell[   10781] = 32'hc123af78;
    ram_cell[   10782] = 32'hde44d2b7;
    ram_cell[   10783] = 32'h8d12fec5;
    ram_cell[   10784] = 32'h09319889;
    ram_cell[   10785] = 32'h9980b5c2;
    ram_cell[   10786] = 32'h4b21ea74;
    ram_cell[   10787] = 32'h9aa6fd02;
    ram_cell[   10788] = 32'h7dbb4e0d;
    ram_cell[   10789] = 32'h6589c222;
    ram_cell[   10790] = 32'hc3ef889f;
    ram_cell[   10791] = 32'ha4aaab88;
    ram_cell[   10792] = 32'hb239c478;
    ram_cell[   10793] = 32'h8f83ec52;
    ram_cell[   10794] = 32'hfb31b2da;
    ram_cell[   10795] = 32'he68f1764;
    ram_cell[   10796] = 32'h064b5419;
    ram_cell[   10797] = 32'hb6ab9abe;
    ram_cell[   10798] = 32'hc36d864a;
    ram_cell[   10799] = 32'h9b52cabe;
    ram_cell[   10800] = 32'h3a07db79;
    ram_cell[   10801] = 32'h8cafc517;
    ram_cell[   10802] = 32'ha1d3a712;
    ram_cell[   10803] = 32'hd3e68637;
    ram_cell[   10804] = 32'hb06df3d4;
    ram_cell[   10805] = 32'hb39f5c96;
    ram_cell[   10806] = 32'hfcfd9b12;
    ram_cell[   10807] = 32'haeda0660;
    ram_cell[   10808] = 32'h42fbbcbc;
    ram_cell[   10809] = 32'h9b48581f;
    ram_cell[   10810] = 32'h21f253ef;
    ram_cell[   10811] = 32'h73ebce0f;
    ram_cell[   10812] = 32'hac6ae374;
    ram_cell[   10813] = 32'h6149ade1;
    ram_cell[   10814] = 32'h4ca747bc;
    ram_cell[   10815] = 32'h55dc1002;
    ram_cell[   10816] = 32'h8ece2af7;
    ram_cell[   10817] = 32'hc9e80abf;
    ram_cell[   10818] = 32'hd5fc09b7;
    ram_cell[   10819] = 32'h1e3390cc;
    ram_cell[   10820] = 32'hc8ac27a3;
    ram_cell[   10821] = 32'h23fb8a80;
    ram_cell[   10822] = 32'h3fa2ae5e;
    ram_cell[   10823] = 32'h177a57e0;
    ram_cell[   10824] = 32'h0a56b62d;
    ram_cell[   10825] = 32'h3e02c3d8;
    ram_cell[   10826] = 32'hb8991c10;
    ram_cell[   10827] = 32'h055caf33;
    ram_cell[   10828] = 32'h57ff4963;
    ram_cell[   10829] = 32'h44a0a40a;
    ram_cell[   10830] = 32'h6a784f89;
    ram_cell[   10831] = 32'h04083606;
    ram_cell[   10832] = 32'h950feaf4;
    ram_cell[   10833] = 32'he1210b44;
    ram_cell[   10834] = 32'hcc9007c9;
    ram_cell[   10835] = 32'h7b7d7f29;
    ram_cell[   10836] = 32'hdde46af7;
    ram_cell[   10837] = 32'h96b21fd2;
    ram_cell[   10838] = 32'h8f8601f5;
    ram_cell[   10839] = 32'h7c5f9cac;
    ram_cell[   10840] = 32'h7fe4cd3c;
    ram_cell[   10841] = 32'hc02323b1;
    ram_cell[   10842] = 32'h7254fde9;
    ram_cell[   10843] = 32'h0d1748e5;
    ram_cell[   10844] = 32'h97786776;
    ram_cell[   10845] = 32'h0a1193bc;
    ram_cell[   10846] = 32'h554ceb4b;
    ram_cell[   10847] = 32'hf8f42ccd;
    ram_cell[   10848] = 32'h1f7e8284;
    ram_cell[   10849] = 32'h4ae29856;
    ram_cell[   10850] = 32'h443624a6;
    ram_cell[   10851] = 32'hbc51f45c;
    ram_cell[   10852] = 32'hbf770145;
    ram_cell[   10853] = 32'ha9a92de0;
    ram_cell[   10854] = 32'h8a796399;
    ram_cell[   10855] = 32'h63e3412b;
    ram_cell[   10856] = 32'h57ea6d4d;
    ram_cell[   10857] = 32'he1d0518f;
    ram_cell[   10858] = 32'h41a31304;
    ram_cell[   10859] = 32'h86d945fc;
    ram_cell[   10860] = 32'heb0a03e4;
    ram_cell[   10861] = 32'he4f586a4;
    ram_cell[   10862] = 32'h47a6b86a;
    ram_cell[   10863] = 32'he6276cde;
    ram_cell[   10864] = 32'hd825b926;
    ram_cell[   10865] = 32'ha3e9115c;
    ram_cell[   10866] = 32'h6491dc1b;
    ram_cell[   10867] = 32'h6a5dcd9a;
    ram_cell[   10868] = 32'h936b51a4;
    ram_cell[   10869] = 32'hc45e1549;
    ram_cell[   10870] = 32'hffd6bcd4;
    ram_cell[   10871] = 32'hfb3d7c64;
    ram_cell[   10872] = 32'hc5268e5d;
    ram_cell[   10873] = 32'he35888ac;
    ram_cell[   10874] = 32'hd99df507;
    ram_cell[   10875] = 32'h37ab7dec;
    ram_cell[   10876] = 32'h968d9ab0;
    ram_cell[   10877] = 32'h8826b83a;
    ram_cell[   10878] = 32'hc834a338;
    ram_cell[   10879] = 32'haf9241a7;
    ram_cell[   10880] = 32'h256057cb;
    ram_cell[   10881] = 32'ha5568dc8;
    ram_cell[   10882] = 32'h9893f29a;
    ram_cell[   10883] = 32'h791cc2a2;
    ram_cell[   10884] = 32'h90a18f04;
    ram_cell[   10885] = 32'hbc099ed7;
    ram_cell[   10886] = 32'h897687a2;
    ram_cell[   10887] = 32'he96b78fe;
    ram_cell[   10888] = 32'h8eef1ac1;
    ram_cell[   10889] = 32'hf2817038;
    ram_cell[   10890] = 32'h18dac94e;
    ram_cell[   10891] = 32'h4d140933;
    ram_cell[   10892] = 32'h24d6df1b;
    ram_cell[   10893] = 32'hf09b91fd;
    ram_cell[   10894] = 32'hcc740bb9;
    ram_cell[   10895] = 32'hddf612ab;
    ram_cell[   10896] = 32'hb61bc550;
    ram_cell[   10897] = 32'h91db0080;
    ram_cell[   10898] = 32'hb29c5990;
    ram_cell[   10899] = 32'h8c90921f;
    ram_cell[   10900] = 32'h55a3a529;
    ram_cell[   10901] = 32'h81e26baa;
    ram_cell[   10902] = 32'had2e9963;
    ram_cell[   10903] = 32'h7a71e446;
    ram_cell[   10904] = 32'hf37d56f8;
    ram_cell[   10905] = 32'h1e48f5b5;
    ram_cell[   10906] = 32'hf98daa2e;
    ram_cell[   10907] = 32'h150d98db;
    ram_cell[   10908] = 32'h4e2ff15f;
    ram_cell[   10909] = 32'h3e040a65;
    ram_cell[   10910] = 32'hae93eec0;
    ram_cell[   10911] = 32'h7298467a;
    ram_cell[   10912] = 32'hd2eb02ed;
    ram_cell[   10913] = 32'h5e26f5ea;
    ram_cell[   10914] = 32'h021da571;
    ram_cell[   10915] = 32'h3238f1f3;
    ram_cell[   10916] = 32'h9d7db31c;
    ram_cell[   10917] = 32'hef76ee7b;
    ram_cell[   10918] = 32'hec1b95ed;
    ram_cell[   10919] = 32'h46d94429;
    ram_cell[   10920] = 32'h3f099caf;
    ram_cell[   10921] = 32'h3bfdbb47;
    ram_cell[   10922] = 32'h6b5161ca;
    ram_cell[   10923] = 32'hd2dc5c9c;
    ram_cell[   10924] = 32'h8fa12ed3;
    ram_cell[   10925] = 32'hae31b2d4;
    ram_cell[   10926] = 32'hd77890d9;
    ram_cell[   10927] = 32'hdeafba1f;
    ram_cell[   10928] = 32'ha387def7;
    ram_cell[   10929] = 32'h6cd3260c;
    ram_cell[   10930] = 32'hb9770848;
    ram_cell[   10931] = 32'he4e5ae8a;
    ram_cell[   10932] = 32'h95a0617e;
    ram_cell[   10933] = 32'hc086fa63;
    ram_cell[   10934] = 32'h33ef594d;
    ram_cell[   10935] = 32'h61e89091;
    ram_cell[   10936] = 32'h8f55e0b3;
    ram_cell[   10937] = 32'hb5154ca4;
    ram_cell[   10938] = 32'hd12cec88;
    ram_cell[   10939] = 32'h9bf3ddf0;
    ram_cell[   10940] = 32'h7d5ea272;
    ram_cell[   10941] = 32'h9aa5e246;
    ram_cell[   10942] = 32'hb1fa929a;
    ram_cell[   10943] = 32'h5567e531;
    ram_cell[   10944] = 32'h96a3110e;
    ram_cell[   10945] = 32'h8e214c53;
    ram_cell[   10946] = 32'h0f134e59;
    ram_cell[   10947] = 32'hfd41417b;
    ram_cell[   10948] = 32'h3958d70e;
    ram_cell[   10949] = 32'hee3bd98e;
    ram_cell[   10950] = 32'hb46ad93d;
    ram_cell[   10951] = 32'ha1d5f134;
    ram_cell[   10952] = 32'h146124d4;
    ram_cell[   10953] = 32'he66f832f;
    ram_cell[   10954] = 32'h97a549b5;
    ram_cell[   10955] = 32'ha900f28c;
    ram_cell[   10956] = 32'h29fdbe52;
    ram_cell[   10957] = 32'hb21ab6cf;
    ram_cell[   10958] = 32'hcaa245e8;
    ram_cell[   10959] = 32'h0c24b8d5;
    ram_cell[   10960] = 32'h33b92626;
    ram_cell[   10961] = 32'h8b2e549f;
    ram_cell[   10962] = 32'h574c6d3d;
    ram_cell[   10963] = 32'h617f4e43;
    ram_cell[   10964] = 32'h4858c7fe;
    ram_cell[   10965] = 32'h155a144c;
    ram_cell[   10966] = 32'h787cab83;
    ram_cell[   10967] = 32'h69266ba8;
    ram_cell[   10968] = 32'hd46824f7;
    ram_cell[   10969] = 32'h9c340208;
    ram_cell[   10970] = 32'hba92b246;
    ram_cell[   10971] = 32'h68c3de02;
    ram_cell[   10972] = 32'hf20a6c14;
    ram_cell[   10973] = 32'h3d4e00d9;
    ram_cell[   10974] = 32'h48d67667;
    ram_cell[   10975] = 32'hccbc3b0f;
    ram_cell[   10976] = 32'h080b0874;
    ram_cell[   10977] = 32'hd1119d96;
    ram_cell[   10978] = 32'hc8ed853f;
    ram_cell[   10979] = 32'h3dbf66b8;
    ram_cell[   10980] = 32'h68afee39;
    ram_cell[   10981] = 32'h44743566;
    ram_cell[   10982] = 32'h8ebc0ef4;
    ram_cell[   10983] = 32'h29ecf7d6;
    ram_cell[   10984] = 32'hbe8571b6;
    ram_cell[   10985] = 32'h2d81c5c0;
    ram_cell[   10986] = 32'hde730ea4;
    ram_cell[   10987] = 32'h39ab5c79;
    ram_cell[   10988] = 32'h69ffa434;
    ram_cell[   10989] = 32'h8b24d76c;
    ram_cell[   10990] = 32'hf498d1ae;
    ram_cell[   10991] = 32'h22df6e8c;
    ram_cell[   10992] = 32'h88ada6ee;
    ram_cell[   10993] = 32'h5b03eeea;
    ram_cell[   10994] = 32'h25a0de0d;
    ram_cell[   10995] = 32'h2f325f60;
    ram_cell[   10996] = 32'hb8df91ee;
    ram_cell[   10997] = 32'h75e09a20;
    ram_cell[   10998] = 32'ha6e29bb5;
    ram_cell[   10999] = 32'hbce27d65;
    ram_cell[   11000] = 32'h40525772;
    ram_cell[   11001] = 32'h6fcd8d8f;
    ram_cell[   11002] = 32'hebcdd870;
    ram_cell[   11003] = 32'h0457edd6;
    ram_cell[   11004] = 32'hc488583d;
    ram_cell[   11005] = 32'hc22e6d63;
    ram_cell[   11006] = 32'h7c9e5d00;
    ram_cell[   11007] = 32'h5051631b;
    ram_cell[   11008] = 32'hba78d6e3;
    ram_cell[   11009] = 32'h78e3448c;
    ram_cell[   11010] = 32'hcd61d75c;
    ram_cell[   11011] = 32'h661a5425;
    ram_cell[   11012] = 32'h5ed2fc66;
    ram_cell[   11013] = 32'h0d0d5fb2;
    ram_cell[   11014] = 32'h823ac9b6;
    ram_cell[   11015] = 32'h09e716f9;
    ram_cell[   11016] = 32'hb119a957;
    ram_cell[   11017] = 32'h8a0d570d;
    ram_cell[   11018] = 32'h76699289;
    ram_cell[   11019] = 32'hefd9b79b;
    ram_cell[   11020] = 32'h77d3d417;
    ram_cell[   11021] = 32'h6e44d654;
    ram_cell[   11022] = 32'h054990af;
    ram_cell[   11023] = 32'h1ba0b687;
    ram_cell[   11024] = 32'h002bf4d0;
    ram_cell[   11025] = 32'hd84de5ee;
    ram_cell[   11026] = 32'h5ff17399;
    ram_cell[   11027] = 32'hf512c9a2;
    ram_cell[   11028] = 32'h5f642248;
    ram_cell[   11029] = 32'h16f80c38;
    ram_cell[   11030] = 32'h3da4566d;
    ram_cell[   11031] = 32'hbc0d6dc7;
    ram_cell[   11032] = 32'hab1d7b77;
    ram_cell[   11033] = 32'hb4626add;
    ram_cell[   11034] = 32'h5c5b1514;
    ram_cell[   11035] = 32'h203f8c3c;
    ram_cell[   11036] = 32'he5c638a0;
    ram_cell[   11037] = 32'h0e796f06;
    ram_cell[   11038] = 32'h4b9e7c74;
    ram_cell[   11039] = 32'h66cb8239;
    ram_cell[   11040] = 32'h7ee30fa7;
    ram_cell[   11041] = 32'hc2498484;
    ram_cell[   11042] = 32'hbbdcd2bc;
    ram_cell[   11043] = 32'h6e7794b8;
    ram_cell[   11044] = 32'hbe58bd5b;
    ram_cell[   11045] = 32'h0feb9f57;
    ram_cell[   11046] = 32'hf0270957;
    ram_cell[   11047] = 32'h4ca17963;
    ram_cell[   11048] = 32'hd0273be6;
    ram_cell[   11049] = 32'hca19617d;
    ram_cell[   11050] = 32'h6521f2be;
    ram_cell[   11051] = 32'h238e9d73;
    ram_cell[   11052] = 32'h293cb625;
    ram_cell[   11053] = 32'h164d21d3;
    ram_cell[   11054] = 32'h3746d0af;
    ram_cell[   11055] = 32'h9c89ac3b;
    ram_cell[   11056] = 32'h94459b88;
    ram_cell[   11057] = 32'h73b0a10f;
    ram_cell[   11058] = 32'h9c4924e6;
    ram_cell[   11059] = 32'h784dcc27;
    ram_cell[   11060] = 32'hc0990430;
    ram_cell[   11061] = 32'h3ca11a02;
    ram_cell[   11062] = 32'h3f2370af;
    ram_cell[   11063] = 32'h7763ca1b;
    ram_cell[   11064] = 32'hc91cd1ad;
    ram_cell[   11065] = 32'h40fc4836;
    ram_cell[   11066] = 32'hd9a937de;
    ram_cell[   11067] = 32'hbf3dd9a6;
    ram_cell[   11068] = 32'h45013b6b;
    ram_cell[   11069] = 32'h1139c5fc;
    ram_cell[   11070] = 32'h0c8e4278;
    ram_cell[   11071] = 32'h0a46bc02;
    ram_cell[   11072] = 32'h69547778;
    ram_cell[   11073] = 32'h58ac2ec3;
    ram_cell[   11074] = 32'h5c7aba49;
    ram_cell[   11075] = 32'hfda82b31;
    ram_cell[   11076] = 32'h26ffccf7;
    ram_cell[   11077] = 32'hf9617392;
    ram_cell[   11078] = 32'hca9d5835;
    ram_cell[   11079] = 32'hb41a8b76;
    ram_cell[   11080] = 32'h8fe1747c;
    ram_cell[   11081] = 32'h09e21a28;
    ram_cell[   11082] = 32'h4f9c3d48;
    ram_cell[   11083] = 32'h0658d266;
    ram_cell[   11084] = 32'h82b99e23;
    ram_cell[   11085] = 32'h1bae8d05;
    ram_cell[   11086] = 32'hf4020588;
    ram_cell[   11087] = 32'h33078bf9;
    ram_cell[   11088] = 32'h2ee3226d;
    ram_cell[   11089] = 32'hd00b51c5;
    ram_cell[   11090] = 32'h9c980b4e;
    ram_cell[   11091] = 32'h40580347;
    ram_cell[   11092] = 32'haf08843b;
    ram_cell[   11093] = 32'hd9c0c47a;
    ram_cell[   11094] = 32'h8b26370c;
    ram_cell[   11095] = 32'hc73931a4;
    ram_cell[   11096] = 32'hf3c8ac21;
    ram_cell[   11097] = 32'h283267d3;
    ram_cell[   11098] = 32'he31e369d;
    ram_cell[   11099] = 32'h9b5e311c;
    ram_cell[   11100] = 32'h63c47c3a;
    ram_cell[   11101] = 32'h28a69107;
    ram_cell[   11102] = 32'hd861bc95;
    ram_cell[   11103] = 32'h97d107b4;
    ram_cell[   11104] = 32'hfe146dd0;
    ram_cell[   11105] = 32'h8986749a;
    ram_cell[   11106] = 32'hf3dfee64;
    ram_cell[   11107] = 32'hefb89e64;
    ram_cell[   11108] = 32'hbc579bfc;
    ram_cell[   11109] = 32'h8aac613d;
    ram_cell[   11110] = 32'h4d975783;
    ram_cell[   11111] = 32'hc1c17919;
    ram_cell[   11112] = 32'h269cc4da;
    ram_cell[   11113] = 32'h0621a929;
    ram_cell[   11114] = 32'h27d489c3;
    ram_cell[   11115] = 32'h595d2bde;
    ram_cell[   11116] = 32'h37faf8d9;
    ram_cell[   11117] = 32'h92d04e77;
    ram_cell[   11118] = 32'he1c44c60;
    ram_cell[   11119] = 32'h70d23b86;
    ram_cell[   11120] = 32'h8e2ba6c6;
    ram_cell[   11121] = 32'hbbbfe109;
    ram_cell[   11122] = 32'h7edd2e89;
    ram_cell[   11123] = 32'h0bdafdb3;
    ram_cell[   11124] = 32'h4465fad2;
    ram_cell[   11125] = 32'h2687c977;
    ram_cell[   11126] = 32'h1af036db;
    ram_cell[   11127] = 32'hfd8be502;
    ram_cell[   11128] = 32'hf8a9c512;
    ram_cell[   11129] = 32'h0efd93a1;
    ram_cell[   11130] = 32'hd52e7ea0;
    ram_cell[   11131] = 32'h7cee786a;
    ram_cell[   11132] = 32'hf2a046c1;
    ram_cell[   11133] = 32'h2224408e;
    ram_cell[   11134] = 32'h11481917;
    ram_cell[   11135] = 32'h1c8cdd2e;
    ram_cell[   11136] = 32'h9d351b9a;
    ram_cell[   11137] = 32'h93fc921e;
    ram_cell[   11138] = 32'h1376b025;
    ram_cell[   11139] = 32'he01acfee;
    ram_cell[   11140] = 32'h4dc4e5a0;
    ram_cell[   11141] = 32'h26678b96;
    ram_cell[   11142] = 32'hf4f2a0b5;
    ram_cell[   11143] = 32'h16b3f404;
    ram_cell[   11144] = 32'h3ca08f5d;
    ram_cell[   11145] = 32'h5a3d5c8d;
    ram_cell[   11146] = 32'h24678166;
    ram_cell[   11147] = 32'hd5752346;
    ram_cell[   11148] = 32'h2a24bcf8;
    ram_cell[   11149] = 32'h6985e9b1;
    ram_cell[   11150] = 32'h078ab2f5;
    ram_cell[   11151] = 32'h8d85e8e6;
    ram_cell[   11152] = 32'h28e860bd;
    ram_cell[   11153] = 32'hff8cacdb;
    ram_cell[   11154] = 32'hc880a008;
    ram_cell[   11155] = 32'h21289983;
    ram_cell[   11156] = 32'h9e37df7c;
    ram_cell[   11157] = 32'hb15dfffe;
    ram_cell[   11158] = 32'hcf47cc8f;
    ram_cell[   11159] = 32'h804e18ec;
    ram_cell[   11160] = 32'h6891ee8b;
    ram_cell[   11161] = 32'h62100815;
    ram_cell[   11162] = 32'h2577ef19;
    ram_cell[   11163] = 32'h5835926c;
    ram_cell[   11164] = 32'hfa274c10;
    ram_cell[   11165] = 32'h0dbfd898;
    ram_cell[   11166] = 32'h188b5149;
    ram_cell[   11167] = 32'h97a76e11;
    ram_cell[   11168] = 32'h8aa77c87;
    ram_cell[   11169] = 32'hfef0f876;
    ram_cell[   11170] = 32'h3267f60d;
    ram_cell[   11171] = 32'h64f4a14f;
    ram_cell[   11172] = 32'h03ed9a12;
    ram_cell[   11173] = 32'hd34bb50d;
    ram_cell[   11174] = 32'h6ae7c0c3;
    ram_cell[   11175] = 32'h04a6d9df;
    ram_cell[   11176] = 32'h76201996;
    ram_cell[   11177] = 32'hc4859cf3;
    ram_cell[   11178] = 32'h65aff172;
    ram_cell[   11179] = 32'h568c0af2;
    ram_cell[   11180] = 32'h30fd089b;
    ram_cell[   11181] = 32'h6b279275;
    ram_cell[   11182] = 32'h22c54b07;
    ram_cell[   11183] = 32'hfd855979;
    ram_cell[   11184] = 32'ha54851c3;
    ram_cell[   11185] = 32'h4c3a9c05;
    ram_cell[   11186] = 32'h8b87bc0a;
    ram_cell[   11187] = 32'h834bb7a9;
    ram_cell[   11188] = 32'hc223b4e8;
    ram_cell[   11189] = 32'h0fc01444;
    ram_cell[   11190] = 32'h67c00c93;
    ram_cell[   11191] = 32'h99ea264c;
    ram_cell[   11192] = 32'h1a373b5d;
    ram_cell[   11193] = 32'h00ac7c15;
    ram_cell[   11194] = 32'h5fdd4d45;
    ram_cell[   11195] = 32'hdde8e627;
    ram_cell[   11196] = 32'h7c1577f1;
    ram_cell[   11197] = 32'hfb428447;
    ram_cell[   11198] = 32'h587101c2;
    ram_cell[   11199] = 32'h583fff43;
    ram_cell[   11200] = 32'hfdb09cc1;
    ram_cell[   11201] = 32'h1140f6ee;
    ram_cell[   11202] = 32'hf90dfa15;
    ram_cell[   11203] = 32'h48cb4f3d;
    ram_cell[   11204] = 32'hb3a15ab5;
    ram_cell[   11205] = 32'hcc7ed312;
    ram_cell[   11206] = 32'h11399d8b;
    ram_cell[   11207] = 32'h2fedb43a;
    ram_cell[   11208] = 32'he083f10c;
    ram_cell[   11209] = 32'hf377b1fd;
    ram_cell[   11210] = 32'h0674d94f;
    ram_cell[   11211] = 32'h72f3bd23;
    ram_cell[   11212] = 32'h42cc403e;
    ram_cell[   11213] = 32'h6eca819c;
    ram_cell[   11214] = 32'hf9911d92;
    ram_cell[   11215] = 32'h30036a0d;
    ram_cell[   11216] = 32'hcd07b397;
    ram_cell[   11217] = 32'hd0a82324;
    ram_cell[   11218] = 32'h58146702;
    ram_cell[   11219] = 32'h643fef11;
    ram_cell[   11220] = 32'h0ca66ac6;
    ram_cell[   11221] = 32'h6703f1b9;
    ram_cell[   11222] = 32'h92c51d88;
    ram_cell[   11223] = 32'hf67e2936;
    ram_cell[   11224] = 32'hc66222ef;
    ram_cell[   11225] = 32'hcc32d35f;
    ram_cell[   11226] = 32'h3e604118;
    ram_cell[   11227] = 32'h04527f8c;
    ram_cell[   11228] = 32'hc65261f3;
    ram_cell[   11229] = 32'h82b4d8c9;
    ram_cell[   11230] = 32'h62e57d3c;
    ram_cell[   11231] = 32'h8866bd34;
    ram_cell[   11232] = 32'h6486670b;
    ram_cell[   11233] = 32'hf30d310e;
    ram_cell[   11234] = 32'h9d2bd732;
    ram_cell[   11235] = 32'h0dc9d271;
    ram_cell[   11236] = 32'h590a81cc;
    ram_cell[   11237] = 32'hd1534223;
    ram_cell[   11238] = 32'h9b4bf6cf;
    ram_cell[   11239] = 32'h71b90a00;
    ram_cell[   11240] = 32'h33c1400c;
    ram_cell[   11241] = 32'h588f6460;
    ram_cell[   11242] = 32'h7ceee014;
    ram_cell[   11243] = 32'h41ddf83b;
    ram_cell[   11244] = 32'h98b31449;
    ram_cell[   11245] = 32'hd50e04ec;
    ram_cell[   11246] = 32'hcd01b4b4;
    ram_cell[   11247] = 32'hdbb8adb6;
    ram_cell[   11248] = 32'h35cec900;
    ram_cell[   11249] = 32'hb1e2fdb3;
    ram_cell[   11250] = 32'h45a6a8f3;
    ram_cell[   11251] = 32'h7bf411ca;
    ram_cell[   11252] = 32'hc5dd7565;
    ram_cell[   11253] = 32'hd4e18862;
    ram_cell[   11254] = 32'h88259a5d;
    ram_cell[   11255] = 32'h8bad33bb;
    ram_cell[   11256] = 32'h4db75713;
    ram_cell[   11257] = 32'h7baa0e1e;
    ram_cell[   11258] = 32'h30c3dae3;
    ram_cell[   11259] = 32'h7230f583;
    ram_cell[   11260] = 32'hfd452fcf;
    ram_cell[   11261] = 32'h6384c271;
    ram_cell[   11262] = 32'h1b8e2ea8;
    ram_cell[   11263] = 32'haa66efc7;
    ram_cell[   11264] = 32'h2eb1460d;
    ram_cell[   11265] = 32'h20ed5ce7;
    ram_cell[   11266] = 32'hd9728c93;
    ram_cell[   11267] = 32'h89212f7b;
    ram_cell[   11268] = 32'h177217a3;
    ram_cell[   11269] = 32'hc20a6fa7;
    ram_cell[   11270] = 32'h8d30ed15;
    ram_cell[   11271] = 32'h0dce35f9;
    ram_cell[   11272] = 32'h2ce364ea;
    ram_cell[   11273] = 32'h046c8f8a;
    ram_cell[   11274] = 32'h81c9dc46;
    ram_cell[   11275] = 32'h1e40cf90;
    ram_cell[   11276] = 32'hcc39ba34;
    ram_cell[   11277] = 32'h912583b3;
    ram_cell[   11278] = 32'hd7e697fa;
    ram_cell[   11279] = 32'hc9ac2db3;
    ram_cell[   11280] = 32'h3b459a32;
    ram_cell[   11281] = 32'h096f8d54;
    ram_cell[   11282] = 32'hddf5dfc8;
    ram_cell[   11283] = 32'h6b0a9c9d;
    ram_cell[   11284] = 32'h32862aa7;
    ram_cell[   11285] = 32'h054204dd;
    ram_cell[   11286] = 32'h15c999be;
    ram_cell[   11287] = 32'h33134490;
    ram_cell[   11288] = 32'h66f78383;
    ram_cell[   11289] = 32'h8da726bc;
    ram_cell[   11290] = 32'he43b68b5;
    ram_cell[   11291] = 32'ha4e775cb;
    ram_cell[   11292] = 32'hbdb1368b;
    ram_cell[   11293] = 32'h8acc02ef;
    ram_cell[   11294] = 32'h84d8c00c;
    ram_cell[   11295] = 32'he84444d5;
    ram_cell[   11296] = 32'h6c652baa;
    ram_cell[   11297] = 32'h57ccebc8;
    ram_cell[   11298] = 32'h5c48bbae;
    ram_cell[   11299] = 32'h34ef4698;
    ram_cell[   11300] = 32'h0a1c8459;
    ram_cell[   11301] = 32'hd7076ab3;
    ram_cell[   11302] = 32'h9b16a97b;
    ram_cell[   11303] = 32'h1c949d97;
    ram_cell[   11304] = 32'h1f561cf7;
    ram_cell[   11305] = 32'h03249973;
    ram_cell[   11306] = 32'hc95d01de;
    ram_cell[   11307] = 32'hff598168;
    ram_cell[   11308] = 32'h4a1e7e0c;
    ram_cell[   11309] = 32'h5c6bf49c;
    ram_cell[   11310] = 32'h8a7c57a4;
    ram_cell[   11311] = 32'ha7439b0b;
    ram_cell[   11312] = 32'h9140f079;
    ram_cell[   11313] = 32'he89c454e;
    ram_cell[   11314] = 32'he26fb0ae;
    ram_cell[   11315] = 32'hbcf19129;
    ram_cell[   11316] = 32'h3f8dd43b;
    ram_cell[   11317] = 32'h96b02251;
    ram_cell[   11318] = 32'ha10f9165;
    ram_cell[   11319] = 32'h56167494;
    ram_cell[   11320] = 32'he21b9f28;
    ram_cell[   11321] = 32'hd64b25f9;
    ram_cell[   11322] = 32'h3fd431a8;
    ram_cell[   11323] = 32'h9449c496;
    ram_cell[   11324] = 32'h49c94730;
    ram_cell[   11325] = 32'hbb1d46f8;
    ram_cell[   11326] = 32'ha7e805e1;
    ram_cell[   11327] = 32'h70748b1f;
    ram_cell[   11328] = 32'hff02dc9f;
    ram_cell[   11329] = 32'heaea0783;
    ram_cell[   11330] = 32'hea538cf6;
    ram_cell[   11331] = 32'h924aef32;
    ram_cell[   11332] = 32'h57ee7ab9;
    ram_cell[   11333] = 32'h46fdc700;
    ram_cell[   11334] = 32'h4c29638e;
    ram_cell[   11335] = 32'ha00fd504;
    ram_cell[   11336] = 32'h71f9f29f;
    ram_cell[   11337] = 32'ha4f832b4;
    ram_cell[   11338] = 32'h1e6e3749;
    ram_cell[   11339] = 32'h919daac0;
    ram_cell[   11340] = 32'ha09f7fcd;
    ram_cell[   11341] = 32'heec74853;
    ram_cell[   11342] = 32'h58d4a93e;
    ram_cell[   11343] = 32'h420d8222;
    ram_cell[   11344] = 32'h9dec043d;
    ram_cell[   11345] = 32'h316557a5;
    ram_cell[   11346] = 32'hf191f3dd;
    ram_cell[   11347] = 32'hff1d7ae4;
    ram_cell[   11348] = 32'h7ff5ad21;
    ram_cell[   11349] = 32'h6c607668;
    ram_cell[   11350] = 32'hbfedb6bd;
    ram_cell[   11351] = 32'h4c5e95f2;
    ram_cell[   11352] = 32'hffcca8b6;
    ram_cell[   11353] = 32'h94f3dabe;
    ram_cell[   11354] = 32'hda6a3f5d;
    ram_cell[   11355] = 32'hb37eb0ef;
    ram_cell[   11356] = 32'hea028b27;
    ram_cell[   11357] = 32'h5e2e0785;
    ram_cell[   11358] = 32'h42328ea4;
    ram_cell[   11359] = 32'hb12b3e27;
    ram_cell[   11360] = 32'hc0b6a0f1;
    ram_cell[   11361] = 32'h9ee803b3;
    ram_cell[   11362] = 32'h8a1bdc7b;
    ram_cell[   11363] = 32'h47cc8788;
    ram_cell[   11364] = 32'hb84debf4;
    ram_cell[   11365] = 32'h6e976de9;
    ram_cell[   11366] = 32'h299eb467;
    ram_cell[   11367] = 32'h43403a00;
    ram_cell[   11368] = 32'h74593ef7;
    ram_cell[   11369] = 32'hb1b56454;
    ram_cell[   11370] = 32'h4000226b;
    ram_cell[   11371] = 32'h7b4d8a46;
    ram_cell[   11372] = 32'he73a770b;
    ram_cell[   11373] = 32'hfb47ffa7;
    ram_cell[   11374] = 32'h3ab33548;
    ram_cell[   11375] = 32'h657708ff;
    ram_cell[   11376] = 32'h6667abaf;
    ram_cell[   11377] = 32'hea036d66;
    ram_cell[   11378] = 32'h9214ca3d;
    ram_cell[   11379] = 32'hc62d5d82;
    ram_cell[   11380] = 32'h95e956b2;
    ram_cell[   11381] = 32'h9082ba18;
    ram_cell[   11382] = 32'hea5d6065;
    ram_cell[   11383] = 32'h71fc3cd4;
    ram_cell[   11384] = 32'h60dcad0a;
    ram_cell[   11385] = 32'h236bc374;
    ram_cell[   11386] = 32'ha9b1b00f;
    ram_cell[   11387] = 32'h091abed3;
    ram_cell[   11388] = 32'h54028f67;
    ram_cell[   11389] = 32'hebb89c86;
    ram_cell[   11390] = 32'h3583a2d6;
    ram_cell[   11391] = 32'h933bb271;
    ram_cell[   11392] = 32'h52d8c1df;
    ram_cell[   11393] = 32'h9fae977a;
    ram_cell[   11394] = 32'hfab296e2;
    ram_cell[   11395] = 32'hbff2067e;
    ram_cell[   11396] = 32'h792bbb22;
    ram_cell[   11397] = 32'hfd03ae1a;
    ram_cell[   11398] = 32'h8f4c0a67;
    ram_cell[   11399] = 32'h7e314879;
    ram_cell[   11400] = 32'h4eb4bc36;
    ram_cell[   11401] = 32'h2379b822;
    ram_cell[   11402] = 32'h446ed127;
    ram_cell[   11403] = 32'h0967db51;
    ram_cell[   11404] = 32'h90e8839b;
    ram_cell[   11405] = 32'hc7fe315c;
    ram_cell[   11406] = 32'h6edb2bd4;
    ram_cell[   11407] = 32'hc7670831;
    ram_cell[   11408] = 32'h96627d04;
    ram_cell[   11409] = 32'h27bb4c41;
    ram_cell[   11410] = 32'h94df9aee;
    ram_cell[   11411] = 32'hbd7970b0;
    ram_cell[   11412] = 32'hd6805875;
    ram_cell[   11413] = 32'h7ad95c53;
    ram_cell[   11414] = 32'h8246f6d0;
    ram_cell[   11415] = 32'hce97f19c;
    ram_cell[   11416] = 32'hc064a187;
    ram_cell[   11417] = 32'hbea5c366;
    ram_cell[   11418] = 32'h63c4c8e5;
    ram_cell[   11419] = 32'h6894e89a;
    ram_cell[   11420] = 32'h20c9b58b;
    ram_cell[   11421] = 32'h300f7daf;
    ram_cell[   11422] = 32'hf3ad113f;
    ram_cell[   11423] = 32'h31d9640d;
    ram_cell[   11424] = 32'h9c4a2474;
    ram_cell[   11425] = 32'h7c61e13c;
    ram_cell[   11426] = 32'haf30d683;
    ram_cell[   11427] = 32'heded6744;
    ram_cell[   11428] = 32'hc86f057a;
    ram_cell[   11429] = 32'h4a2e84b9;
    ram_cell[   11430] = 32'hd8f2b146;
    ram_cell[   11431] = 32'h22166007;
    ram_cell[   11432] = 32'ha3ad4649;
    ram_cell[   11433] = 32'hd98f9dc5;
    ram_cell[   11434] = 32'h78a97da2;
    ram_cell[   11435] = 32'h9b9e1b96;
    ram_cell[   11436] = 32'h229992b4;
    ram_cell[   11437] = 32'he13b17f4;
    ram_cell[   11438] = 32'hc07b5b90;
    ram_cell[   11439] = 32'hecd11bf8;
    ram_cell[   11440] = 32'hbdf850ee;
    ram_cell[   11441] = 32'h78734d67;
    ram_cell[   11442] = 32'hb5f336b0;
    ram_cell[   11443] = 32'h4e78309d;
    ram_cell[   11444] = 32'h608ab48c;
    ram_cell[   11445] = 32'h76770568;
    ram_cell[   11446] = 32'hb88883ce;
    ram_cell[   11447] = 32'h49045782;
    ram_cell[   11448] = 32'h77f24d2d;
    ram_cell[   11449] = 32'hdd6ba5f9;
    ram_cell[   11450] = 32'h0c87b6a0;
    ram_cell[   11451] = 32'h9755a4b1;
    ram_cell[   11452] = 32'hdd4f166e;
    ram_cell[   11453] = 32'h787c8323;
    ram_cell[   11454] = 32'h9da96368;
    ram_cell[   11455] = 32'h6a5a965c;
    ram_cell[   11456] = 32'h35d186ce;
    ram_cell[   11457] = 32'h1a25076b;
    ram_cell[   11458] = 32'hcabf6eee;
    ram_cell[   11459] = 32'h0c6e00b4;
    ram_cell[   11460] = 32'he695f103;
    ram_cell[   11461] = 32'hc48c3cc5;
    ram_cell[   11462] = 32'hf24cf8e8;
    ram_cell[   11463] = 32'h1b437503;
    ram_cell[   11464] = 32'he227b1c8;
    ram_cell[   11465] = 32'hcd68991a;
    ram_cell[   11466] = 32'h835c1697;
    ram_cell[   11467] = 32'ha8d42e28;
    ram_cell[   11468] = 32'h672baa33;
    ram_cell[   11469] = 32'haa598e06;
    ram_cell[   11470] = 32'h39d18e81;
    ram_cell[   11471] = 32'hdcd080fb;
    ram_cell[   11472] = 32'h159bad58;
    ram_cell[   11473] = 32'he4711750;
    ram_cell[   11474] = 32'h27647aa3;
    ram_cell[   11475] = 32'h83aa1dd3;
    ram_cell[   11476] = 32'h8bd01b7d;
    ram_cell[   11477] = 32'ha34d3b8c;
    ram_cell[   11478] = 32'h85775bdd;
    ram_cell[   11479] = 32'hecf5a0a0;
    ram_cell[   11480] = 32'h534e503e;
    ram_cell[   11481] = 32'he2bda942;
    ram_cell[   11482] = 32'h207ce221;
    ram_cell[   11483] = 32'h10d11631;
    ram_cell[   11484] = 32'h39559971;
    ram_cell[   11485] = 32'h32a81122;
    ram_cell[   11486] = 32'hd781e214;
    ram_cell[   11487] = 32'h6a32dcf1;
    ram_cell[   11488] = 32'ha2313094;
    ram_cell[   11489] = 32'h90185131;
    ram_cell[   11490] = 32'h639d9b5f;
    ram_cell[   11491] = 32'ha622082c;
    ram_cell[   11492] = 32'hbe95313c;
    ram_cell[   11493] = 32'hdf8fbb93;
    ram_cell[   11494] = 32'h5b011cef;
    ram_cell[   11495] = 32'h2396e1c2;
    ram_cell[   11496] = 32'hdd84fef3;
    ram_cell[   11497] = 32'h1b9506fb;
    ram_cell[   11498] = 32'h6c410e88;
    ram_cell[   11499] = 32'h2c2fa2a0;
    ram_cell[   11500] = 32'he1875380;
    ram_cell[   11501] = 32'h23db24f6;
    ram_cell[   11502] = 32'hceba122f;
    ram_cell[   11503] = 32'h1c78e5ed;
    ram_cell[   11504] = 32'h81f6371a;
    ram_cell[   11505] = 32'h62b10915;
    ram_cell[   11506] = 32'h381e366b;
    ram_cell[   11507] = 32'habe08807;
    ram_cell[   11508] = 32'h96a670f2;
    ram_cell[   11509] = 32'h48eb21d8;
    ram_cell[   11510] = 32'hc5dcd9f8;
    ram_cell[   11511] = 32'h144a443c;
    ram_cell[   11512] = 32'h75f3b531;
    ram_cell[   11513] = 32'ha67c089b;
    ram_cell[   11514] = 32'h5c8d04fb;
    ram_cell[   11515] = 32'hf6d1e1ba;
    ram_cell[   11516] = 32'h7e72f31c;
    ram_cell[   11517] = 32'h92cdc937;
    ram_cell[   11518] = 32'hf62301fd;
    ram_cell[   11519] = 32'he75e38b9;
    ram_cell[   11520] = 32'h48116046;
    ram_cell[   11521] = 32'h35a74842;
    ram_cell[   11522] = 32'h512ce218;
    ram_cell[   11523] = 32'h0123f6f2;
    ram_cell[   11524] = 32'h8b2d1a3f;
    ram_cell[   11525] = 32'h15624e89;
    ram_cell[   11526] = 32'h157ed996;
    ram_cell[   11527] = 32'hb774b739;
    ram_cell[   11528] = 32'h07021eb3;
    ram_cell[   11529] = 32'h56d407b4;
    ram_cell[   11530] = 32'hf1f1663b;
    ram_cell[   11531] = 32'h6bc3ee6c;
    ram_cell[   11532] = 32'h9d6284eb;
    ram_cell[   11533] = 32'h932fd88a;
    ram_cell[   11534] = 32'ha0615ce9;
    ram_cell[   11535] = 32'h2bcb4323;
    ram_cell[   11536] = 32'hfd578cb6;
    ram_cell[   11537] = 32'hd4232ddf;
    ram_cell[   11538] = 32'hcaa09152;
    ram_cell[   11539] = 32'h9ccfdba2;
    ram_cell[   11540] = 32'h4f8ece7a;
    ram_cell[   11541] = 32'h85a59829;
    ram_cell[   11542] = 32'ha9e637ff;
    ram_cell[   11543] = 32'h37445c58;
    ram_cell[   11544] = 32'h1fc9ca24;
    ram_cell[   11545] = 32'h2cf10b27;
    ram_cell[   11546] = 32'h940cc132;
    ram_cell[   11547] = 32'hcbfce744;
    ram_cell[   11548] = 32'h3a9c377e;
    ram_cell[   11549] = 32'ha2ed03ca;
    ram_cell[   11550] = 32'h815d3162;
    ram_cell[   11551] = 32'h80adaccf;
    ram_cell[   11552] = 32'hbf58bb04;
    ram_cell[   11553] = 32'h4410edff;
    ram_cell[   11554] = 32'h96409694;
    ram_cell[   11555] = 32'h824baed4;
    ram_cell[   11556] = 32'h51ab9734;
    ram_cell[   11557] = 32'h6c42956c;
    ram_cell[   11558] = 32'h829854f4;
    ram_cell[   11559] = 32'h9da6e644;
    ram_cell[   11560] = 32'h24f15ad5;
    ram_cell[   11561] = 32'h48834581;
    ram_cell[   11562] = 32'hbc1cc565;
    ram_cell[   11563] = 32'h0fbe781c;
    ram_cell[   11564] = 32'hf9213f30;
    ram_cell[   11565] = 32'h6f8a59e0;
    ram_cell[   11566] = 32'h2d6951c2;
    ram_cell[   11567] = 32'h54e73507;
    ram_cell[   11568] = 32'h1382d2b9;
    ram_cell[   11569] = 32'h298a0fd7;
    ram_cell[   11570] = 32'h51c9d53d;
    ram_cell[   11571] = 32'he2485d7e;
    ram_cell[   11572] = 32'h19639521;
    ram_cell[   11573] = 32'h00e9543a;
    ram_cell[   11574] = 32'haf3ca207;
    ram_cell[   11575] = 32'h94d40a3a;
    ram_cell[   11576] = 32'hfeee6c22;
    ram_cell[   11577] = 32'h754f60f2;
    ram_cell[   11578] = 32'hbb53ec00;
    ram_cell[   11579] = 32'h2b5214d0;
    ram_cell[   11580] = 32'h2ac9438e;
    ram_cell[   11581] = 32'hdf755525;
    ram_cell[   11582] = 32'h6e77c9a3;
    ram_cell[   11583] = 32'hf250c4c1;
    ram_cell[   11584] = 32'h75f35317;
    ram_cell[   11585] = 32'h254257df;
    ram_cell[   11586] = 32'h1c12b134;
    ram_cell[   11587] = 32'h91ea03f9;
    ram_cell[   11588] = 32'h6427f380;
    ram_cell[   11589] = 32'hdb3fa375;
    ram_cell[   11590] = 32'ha10884ca;
    ram_cell[   11591] = 32'h69d5b56b;
    ram_cell[   11592] = 32'h10fdcc62;
    ram_cell[   11593] = 32'h721490bf;
    ram_cell[   11594] = 32'heb23dd74;
    ram_cell[   11595] = 32'hfa012916;
    ram_cell[   11596] = 32'hf7f7caa0;
    ram_cell[   11597] = 32'hae189172;
    ram_cell[   11598] = 32'h6ae67c75;
    ram_cell[   11599] = 32'h05e66491;
    ram_cell[   11600] = 32'hee5f520b;
    ram_cell[   11601] = 32'h240583ef;
    ram_cell[   11602] = 32'h4425332d;
    ram_cell[   11603] = 32'he1bbf157;
    ram_cell[   11604] = 32'h4806a324;
    ram_cell[   11605] = 32'h4ffce317;
    ram_cell[   11606] = 32'hb5488128;
    ram_cell[   11607] = 32'h95f92379;
    ram_cell[   11608] = 32'hcb723357;
    ram_cell[   11609] = 32'hdab12f89;
    ram_cell[   11610] = 32'h92acca64;
    ram_cell[   11611] = 32'h11af779b;
    ram_cell[   11612] = 32'hb129dcd6;
    ram_cell[   11613] = 32'hd0c51ed9;
    ram_cell[   11614] = 32'h127ffc54;
    ram_cell[   11615] = 32'h04c66380;
    ram_cell[   11616] = 32'hc8a2442e;
    ram_cell[   11617] = 32'h017305cf;
    ram_cell[   11618] = 32'h1d276973;
    ram_cell[   11619] = 32'hb9984578;
    ram_cell[   11620] = 32'hf4612e9f;
    ram_cell[   11621] = 32'hafa5391b;
    ram_cell[   11622] = 32'haef06c50;
    ram_cell[   11623] = 32'h9b903f91;
    ram_cell[   11624] = 32'hcad1f95f;
    ram_cell[   11625] = 32'hf56027a4;
    ram_cell[   11626] = 32'h0abf6ec8;
    ram_cell[   11627] = 32'h8e36d9b8;
    ram_cell[   11628] = 32'h2b3990f0;
    ram_cell[   11629] = 32'h14df553d;
    ram_cell[   11630] = 32'h3f815c45;
    ram_cell[   11631] = 32'h24187d97;
    ram_cell[   11632] = 32'hcd378ee2;
    ram_cell[   11633] = 32'h53e3bbeb;
    ram_cell[   11634] = 32'hea4f6209;
    ram_cell[   11635] = 32'ha181ce82;
    ram_cell[   11636] = 32'h65f73e07;
    ram_cell[   11637] = 32'hf86681b1;
    ram_cell[   11638] = 32'h9e26199b;
    ram_cell[   11639] = 32'h02c3c881;
    ram_cell[   11640] = 32'h387d0023;
    ram_cell[   11641] = 32'h65ca3a4f;
    ram_cell[   11642] = 32'h62214252;
    ram_cell[   11643] = 32'hccd83f9e;
    ram_cell[   11644] = 32'h33d07ec8;
    ram_cell[   11645] = 32'h5eb5e07e;
    ram_cell[   11646] = 32'hb9e3f0d3;
    ram_cell[   11647] = 32'h99d4a688;
    ram_cell[   11648] = 32'hcd232e81;
    ram_cell[   11649] = 32'h14c57414;
    ram_cell[   11650] = 32'h624f53a0;
    ram_cell[   11651] = 32'h591c132e;
    ram_cell[   11652] = 32'he323c13d;
    ram_cell[   11653] = 32'h9450732f;
    ram_cell[   11654] = 32'h0231d648;
    ram_cell[   11655] = 32'h129f1c8b;
    ram_cell[   11656] = 32'h50f40dbd;
    ram_cell[   11657] = 32'h08f76f19;
    ram_cell[   11658] = 32'h711b6725;
    ram_cell[   11659] = 32'hc5d3c13e;
    ram_cell[   11660] = 32'hecbcd935;
    ram_cell[   11661] = 32'h944b2d74;
    ram_cell[   11662] = 32'hc829f4fb;
    ram_cell[   11663] = 32'h1b00044a;
    ram_cell[   11664] = 32'h0445b56b;
    ram_cell[   11665] = 32'hb5cd723d;
    ram_cell[   11666] = 32'h2a1ca997;
    ram_cell[   11667] = 32'hee6881ec;
    ram_cell[   11668] = 32'h075a2635;
    ram_cell[   11669] = 32'h0983e382;
    ram_cell[   11670] = 32'hd315ccdc;
    ram_cell[   11671] = 32'h8577566c;
    ram_cell[   11672] = 32'h5e752433;
    ram_cell[   11673] = 32'h859ee1fe;
    ram_cell[   11674] = 32'he4dfb58a;
    ram_cell[   11675] = 32'ha50e9475;
    ram_cell[   11676] = 32'ha333a42d;
    ram_cell[   11677] = 32'hf6f858b3;
    ram_cell[   11678] = 32'hd0f887e4;
    ram_cell[   11679] = 32'h880fc2cd;
    ram_cell[   11680] = 32'hb5e46248;
    ram_cell[   11681] = 32'he13fe35b;
    ram_cell[   11682] = 32'h4cb9d5b9;
    ram_cell[   11683] = 32'h0c11a03b;
    ram_cell[   11684] = 32'h9aa97eb8;
    ram_cell[   11685] = 32'h465b0104;
    ram_cell[   11686] = 32'he1e04764;
    ram_cell[   11687] = 32'h1f8d5401;
    ram_cell[   11688] = 32'h9c4a049f;
    ram_cell[   11689] = 32'he2c72614;
    ram_cell[   11690] = 32'h05177c16;
    ram_cell[   11691] = 32'h98694850;
    ram_cell[   11692] = 32'hc9651e01;
    ram_cell[   11693] = 32'h26f56fbc;
    ram_cell[   11694] = 32'hab2f45dd;
    ram_cell[   11695] = 32'ha1c432eb;
    ram_cell[   11696] = 32'h684e4819;
    ram_cell[   11697] = 32'hffa0ad14;
    ram_cell[   11698] = 32'ha4fba479;
    ram_cell[   11699] = 32'hee5d758f;
    ram_cell[   11700] = 32'h8b68c910;
    ram_cell[   11701] = 32'hfee7a3e7;
    ram_cell[   11702] = 32'hdc8fc2c1;
    ram_cell[   11703] = 32'h6855aab8;
    ram_cell[   11704] = 32'hbc555b89;
    ram_cell[   11705] = 32'h10be82d0;
    ram_cell[   11706] = 32'hf256c175;
    ram_cell[   11707] = 32'h2b7b5012;
    ram_cell[   11708] = 32'h78d00a30;
    ram_cell[   11709] = 32'h75754a5a;
    ram_cell[   11710] = 32'h0f8986df;
    ram_cell[   11711] = 32'h6eb733b5;
    ram_cell[   11712] = 32'hbf85909b;
    ram_cell[   11713] = 32'hcc231fa6;
    ram_cell[   11714] = 32'h38f425a2;
    ram_cell[   11715] = 32'h9f2a8aa6;
    ram_cell[   11716] = 32'h74ad39bb;
    ram_cell[   11717] = 32'h01a45d93;
    ram_cell[   11718] = 32'h3e4b9ad1;
    ram_cell[   11719] = 32'heee54430;
    ram_cell[   11720] = 32'h1fa121fb;
    ram_cell[   11721] = 32'h149f009c;
    ram_cell[   11722] = 32'hcc633960;
    ram_cell[   11723] = 32'h3593c867;
    ram_cell[   11724] = 32'h6ed4dd96;
    ram_cell[   11725] = 32'h4397d596;
    ram_cell[   11726] = 32'hb76fe027;
    ram_cell[   11727] = 32'h4709a1e2;
    ram_cell[   11728] = 32'hb86fb078;
    ram_cell[   11729] = 32'ha040374d;
    ram_cell[   11730] = 32'hf96583ed;
    ram_cell[   11731] = 32'h3e1950c2;
    ram_cell[   11732] = 32'h958ae777;
    ram_cell[   11733] = 32'h43bc024d;
    ram_cell[   11734] = 32'h2e89a98f;
    ram_cell[   11735] = 32'hd3ae9907;
    ram_cell[   11736] = 32'hf73d1208;
    ram_cell[   11737] = 32'he9fa7f81;
    ram_cell[   11738] = 32'h2782f419;
    ram_cell[   11739] = 32'h039e3b33;
    ram_cell[   11740] = 32'h7df844c2;
    ram_cell[   11741] = 32'ha9709f92;
    ram_cell[   11742] = 32'h93ff5370;
    ram_cell[   11743] = 32'h5750dbd0;
    ram_cell[   11744] = 32'h1c1a1901;
    ram_cell[   11745] = 32'h10e58f71;
    ram_cell[   11746] = 32'h426a78bb;
    ram_cell[   11747] = 32'hb1003cb2;
    ram_cell[   11748] = 32'hb9985faf;
    ram_cell[   11749] = 32'h25841921;
    ram_cell[   11750] = 32'hf73a0948;
    ram_cell[   11751] = 32'h764a0ced;
    ram_cell[   11752] = 32'h34db9e0d;
    ram_cell[   11753] = 32'h281b5a20;
    ram_cell[   11754] = 32'h6e0133a1;
    ram_cell[   11755] = 32'hcaaf2785;
    ram_cell[   11756] = 32'h3c8f9790;
    ram_cell[   11757] = 32'hae3cabc2;
    ram_cell[   11758] = 32'h46ee6d61;
    ram_cell[   11759] = 32'h4696acbc;
    ram_cell[   11760] = 32'haaf40f5d;
    ram_cell[   11761] = 32'he39c76f8;
    ram_cell[   11762] = 32'h0e586050;
    ram_cell[   11763] = 32'ha9e06a10;
    ram_cell[   11764] = 32'h02ceacd9;
    ram_cell[   11765] = 32'h47800b1c;
    ram_cell[   11766] = 32'h4cbd89e6;
    ram_cell[   11767] = 32'h3ed4495e;
    ram_cell[   11768] = 32'h662d7cfb;
    ram_cell[   11769] = 32'h17a4025d;
    ram_cell[   11770] = 32'hb3f1ea6a;
    ram_cell[   11771] = 32'h29d479f9;
    ram_cell[   11772] = 32'hdd6fa647;
    ram_cell[   11773] = 32'hf09ca2c3;
    ram_cell[   11774] = 32'h3e7874ce;
    ram_cell[   11775] = 32'h1df24fe7;
    ram_cell[   11776] = 32'haec7bc2c;
    ram_cell[   11777] = 32'h6e381d37;
    ram_cell[   11778] = 32'h2d5942c1;
    ram_cell[   11779] = 32'h4ea50b20;
    ram_cell[   11780] = 32'hcd0acc3a;
    ram_cell[   11781] = 32'hc5c768a5;
    ram_cell[   11782] = 32'h2f8e92eb;
    ram_cell[   11783] = 32'heb0db1a9;
    ram_cell[   11784] = 32'hf72e35b3;
    ram_cell[   11785] = 32'h7be01e40;
    ram_cell[   11786] = 32'h99bc98f5;
    ram_cell[   11787] = 32'h17cc0cfb;
    ram_cell[   11788] = 32'hf49da236;
    ram_cell[   11789] = 32'he3c31a8c;
    ram_cell[   11790] = 32'h2ac801c7;
    ram_cell[   11791] = 32'h9cf97244;
    ram_cell[   11792] = 32'h67cc27cf;
    ram_cell[   11793] = 32'hcaf2df9d;
    ram_cell[   11794] = 32'heda0b1a5;
    ram_cell[   11795] = 32'ha2b445dc;
    ram_cell[   11796] = 32'h593b0bdf;
    ram_cell[   11797] = 32'h01ea54b5;
    ram_cell[   11798] = 32'h4137c4c5;
    ram_cell[   11799] = 32'h3d5c2717;
    ram_cell[   11800] = 32'hdea76d04;
    ram_cell[   11801] = 32'h49a32a25;
    ram_cell[   11802] = 32'he347d71a;
    ram_cell[   11803] = 32'h4343fa57;
    ram_cell[   11804] = 32'hfb875d23;
    ram_cell[   11805] = 32'h93749fde;
    ram_cell[   11806] = 32'h2fd2b33c;
    ram_cell[   11807] = 32'hfceb4c83;
    ram_cell[   11808] = 32'h9cefa25a;
    ram_cell[   11809] = 32'h77d94e2f;
    ram_cell[   11810] = 32'h74bc0ea2;
    ram_cell[   11811] = 32'hb99290d6;
    ram_cell[   11812] = 32'h5797bce5;
    ram_cell[   11813] = 32'had8e9dc0;
    ram_cell[   11814] = 32'h43eb318d;
    ram_cell[   11815] = 32'h8835dcc6;
    ram_cell[   11816] = 32'h9d12057c;
    ram_cell[   11817] = 32'h2a4750b8;
    ram_cell[   11818] = 32'h4a861de8;
    ram_cell[   11819] = 32'h87a1d946;
    ram_cell[   11820] = 32'h14cd9f2c;
    ram_cell[   11821] = 32'hac82ef9f;
    ram_cell[   11822] = 32'h32ea44ee;
    ram_cell[   11823] = 32'he1aef7db;
    ram_cell[   11824] = 32'hcca72065;
    ram_cell[   11825] = 32'hd40103fa;
    ram_cell[   11826] = 32'h82a8dd5f;
    ram_cell[   11827] = 32'h5ade2caf;
    ram_cell[   11828] = 32'h60b7b0fe;
    ram_cell[   11829] = 32'h420481eb;
    ram_cell[   11830] = 32'h1013a295;
    ram_cell[   11831] = 32'hfc128f54;
    ram_cell[   11832] = 32'hc7526dea;
    ram_cell[   11833] = 32'h0b27f41a;
    ram_cell[   11834] = 32'hc6839384;
    ram_cell[   11835] = 32'hb0cac8fb;
    ram_cell[   11836] = 32'h5cecd5a2;
    ram_cell[   11837] = 32'h3c85c72f;
    ram_cell[   11838] = 32'hd83f7116;
    ram_cell[   11839] = 32'h69dbea73;
    ram_cell[   11840] = 32'h8a6d8b41;
    ram_cell[   11841] = 32'hd6857da3;
    ram_cell[   11842] = 32'h6af4dfd5;
    ram_cell[   11843] = 32'ha56fa8e1;
    ram_cell[   11844] = 32'hfdb8832b;
    ram_cell[   11845] = 32'h39285160;
    ram_cell[   11846] = 32'h82f1c03c;
    ram_cell[   11847] = 32'ha0141c56;
    ram_cell[   11848] = 32'hd9f37697;
    ram_cell[   11849] = 32'h9a58b8ae;
    ram_cell[   11850] = 32'ha549f91c;
    ram_cell[   11851] = 32'hc6ba8d88;
    ram_cell[   11852] = 32'h7e84d630;
    ram_cell[   11853] = 32'hf0239773;
    ram_cell[   11854] = 32'h152a760c;
    ram_cell[   11855] = 32'h124e1279;
    ram_cell[   11856] = 32'h6e5b47d7;
    ram_cell[   11857] = 32'hb1f034d9;
    ram_cell[   11858] = 32'h54b07399;
    ram_cell[   11859] = 32'h7a2e59e2;
    ram_cell[   11860] = 32'h08d33d78;
    ram_cell[   11861] = 32'h9c1443ab;
    ram_cell[   11862] = 32'haec6489d;
    ram_cell[   11863] = 32'h4709f55b;
    ram_cell[   11864] = 32'hafef135e;
    ram_cell[   11865] = 32'h5abd2dad;
    ram_cell[   11866] = 32'h1b6cf74c;
    ram_cell[   11867] = 32'hd9371c66;
    ram_cell[   11868] = 32'h9ee7b23a;
    ram_cell[   11869] = 32'hb6f2f29b;
    ram_cell[   11870] = 32'hb7da6baa;
    ram_cell[   11871] = 32'hde830ae6;
    ram_cell[   11872] = 32'hae250db1;
    ram_cell[   11873] = 32'h79d5b6f2;
    ram_cell[   11874] = 32'h760384ca;
    ram_cell[   11875] = 32'h2b5e6f28;
    ram_cell[   11876] = 32'h8904ec75;
    ram_cell[   11877] = 32'h5df379d2;
    ram_cell[   11878] = 32'h1e4e4306;
    ram_cell[   11879] = 32'h15ab3c77;
    ram_cell[   11880] = 32'h7d2149f9;
    ram_cell[   11881] = 32'h7e466618;
    ram_cell[   11882] = 32'h510b5bf2;
    ram_cell[   11883] = 32'hda95f7a5;
    ram_cell[   11884] = 32'he68a1c12;
    ram_cell[   11885] = 32'ha30e021e;
    ram_cell[   11886] = 32'h05734349;
    ram_cell[   11887] = 32'ha11ef562;
    ram_cell[   11888] = 32'h7e992b06;
    ram_cell[   11889] = 32'h47aee649;
    ram_cell[   11890] = 32'h40247a78;
    ram_cell[   11891] = 32'ha61c468e;
    ram_cell[   11892] = 32'hd93566bb;
    ram_cell[   11893] = 32'h371d24fa;
    ram_cell[   11894] = 32'hbbb54f39;
    ram_cell[   11895] = 32'hb559c359;
    ram_cell[   11896] = 32'h86c8d75d;
    ram_cell[   11897] = 32'hb4db7ed9;
    ram_cell[   11898] = 32'h7b2f9e71;
    ram_cell[   11899] = 32'hdb8dcd33;
    ram_cell[   11900] = 32'h9dadb445;
    ram_cell[   11901] = 32'h510503c5;
    ram_cell[   11902] = 32'h373f079c;
    ram_cell[   11903] = 32'h7cc73954;
    ram_cell[   11904] = 32'hce0b757f;
    ram_cell[   11905] = 32'h78da8e57;
    ram_cell[   11906] = 32'h6042bc36;
    ram_cell[   11907] = 32'h0400eb6e;
    ram_cell[   11908] = 32'h68322620;
    ram_cell[   11909] = 32'h023f77c5;
    ram_cell[   11910] = 32'h9a01d812;
    ram_cell[   11911] = 32'ha8549447;
    ram_cell[   11912] = 32'hd9b92f87;
    ram_cell[   11913] = 32'h72af3824;
    ram_cell[   11914] = 32'hb84862ee;
    ram_cell[   11915] = 32'hd720616a;
    ram_cell[   11916] = 32'h3881d951;
    ram_cell[   11917] = 32'hf8590da0;
    ram_cell[   11918] = 32'h46fc32c4;
    ram_cell[   11919] = 32'hd1364514;
    ram_cell[   11920] = 32'h2a4c92d5;
    ram_cell[   11921] = 32'h33cb2ef9;
    ram_cell[   11922] = 32'hac5dcb55;
    ram_cell[   11923] = 32'h401fb36e;
    ram_cell[   11924] = 32'h1d36fe7e;
    ram_cell[   11925] = 32'hb72463ff;
    ram_cell[   11926] = 32'hca2151b4;
    ram_cell[   11927] = 32'h6a86d33b;
    ram_cell[   11928] = 32'h8969cde6;
    ram_cell[   11929] = 32'hcb4c3b47;
    ram_cell[   11930] = 32'h6e763d6f;
    ram_cell[   11931] = 32'hd124635e;
    ram_cell[   11932] = 32'h11a74a39;
    ram_cell[   11933] = 32'h535be16c;
    ram_cell[   11934] = 32'h0e84f670;
    ram_cell[   11935] = 32'h42283fe2;
    ram_cell[   11936] = 32'h07bc5068;
    ram_cell[   11937] = 32'h9dc504cb;
    ram_cell[   11938] = 32'hf9b8ee55;
    ram_cell[   11939] = 32'h22e8579d;
    ram_cell[   11940] = 32'hbb8a76a1;
    ram_cell[   11941] = 32'hfbf8d338;
    ram_cell[   11942] = 32'hf45687ad;
    ram_cell[   11943] = 32'h8e5d0a08;
    ram_cell[   11944] = 32'h9b096e6c;
    ram_cell[   11945] = 32'h583e60a4;
    ram_cell[   11946] = 32'h3da7e34a;
    ram_cell[   11947] = 32'hdb4c6915;
    ram_cell[   11948] = 32'he227dc39;
    ram_cell[   11949] = 32'h4f8ff186;
    ram_cell[   11950] = 32'h9d9c1f0e;
    ram_cell[   11951] = 32'h5e39aaa7;
    ram_cell[   11952] = 32'h90ec2b29;
    ram_cell[   11953] = 32'hd5e1a2bf;
    ram_cell[   11954] = 32'h0a25d13a;
    ram_cell[   11955] = 32'h67df2511;
    ram_cell[   11956] = 32'hde1df61a;
    ram_cell[   11957] = 32'h1b44e21a;
    ram_cell[   11958] = 32'hfc26c15e;
    ram_cell[   11959] = 32'h7f6b47fa;
    ram_cell[   11960] = 32'h7bea9b8c;
    ram_cell[   11961] = 32'h739ba0ad;
    ram_cell[   11962] = 32'ha6d737de;
    ram_cell[   11963] = 32'h76e59682;
    ram_cell[   11964] = 32'h9bbca10d;
    ram_cell[   11965] = 32'h05d76725;
    ram_cell[   11966] = 32'h7f8dfc55;
    ram_cell[   11967] = 32'h432aeec6;
    ram_cell[   11968] = 32'h7f627213;
    ram_cell[   11969] = 32'hd4814ef1;
    ram_cell[   11970] = 32'h837bf8f2;
    ram_cell[   11971] = 32'h5d1fb240;
    ram_cell[   11972] = 32'hc9907082;
    ram_cell[   11973] = 32'haabd8533;
    ram_cell[   11974] = 32'h30556874;
    ram_cell[   11975] = 32'h233be74f;
    ram_cell[   11976] = 32'h59610f64;
    ram_cell[   11977] = 32'h97d76cd2;
    ram_cell[   11978] = 32'hcc122f5b;
    ram_cell[   11979] = 32'haaeb98bf;
    ram_cell[   11980] = 32'hb4a6d954;
    ram_cell[   11981] = 32'h0cf14edd;
    ram_cell[   11982] = 32'h4181846c;
    ram_cell[   11983] = 32'h71ef37af;
    ram_cell[   11984] = 32'h941a05c1;
    ram_cell[   11985] = 32'h7e8aeb72;
    ram_cell[   11986] = 32'h0e51d278;
    ram_cell[   11987] = 32'h591db654;
    ram_cell[   11988] = 32'hba27fec5;
    ram_cell[   11989] = 32'h422da86e;
    ram_cell[   11990] = 32'h188cb84d;
    ram_cell[   11991] = 32'h9be429df;
    ram_cell[   11992] = 32'h7cbb2bad;
    ram_cell[   11993] = 32'h4a99f154;
    ram_cell[   11994] = 32'h097cf5f2;
    ram_cell[   11995] = 32'h0c8efc50;
    ram_cell[   11996] = 32'h435d766c;
    ram_cell[   11997] = 32'h60332ac6;
    ram_cell[   11998] = 32'h51ceec0d;
    ram_cell[   11999] = 32'hadf51a4b;
    ram_cell[   12000] = 32'h9e284e8c;
    ram_cell[   12001] = 32'hcfadb109;
    ram_cell[   12002] = 32'h5a6d15cb;
    ram_cell[   12003] = 32'hc02dd84c;
    ram_cell[   12004] = 32'haae4ce33;
    ram_cell[   12005] = 32'h2983838a;
    ram_cell[   12006] = 32'hcfc27444;
    ram_cell[   12007] = 32'h3bcf881d;
    ram_cell[   12008] = 32'h2d2df77b;
    ram_cell[   12009] = 32'h54edafc3;
    ram_cell[   12010] = 32'hd99a8338;
    ram_cell[   12011] = 32'h653f4472;
    ram_cell[   12012] = 32'hec9420c5;
    ram_cell[   12013] = 32'h88be5889;
    ram_cell[   12014] = 32'h8267f8e9;
    ram_cell[   12015] = 32'hd8336770;
    ram_cell[   12016] = 32'hf8b11aea;
    ram_cell[   12017] = 32'ha79b0e22;
    ram_cell[   12018] = 32'he4549a5a;
    ram_cell[   12019] = 32'h715e531e;
    ram_cell[   12020] = 32'hb95e2b18;
    ram_cell[   12021] = 32'ha49f53ed;
    ram_cell[   12022] = 32'hcdad1e17;
    ram_cell[   12023] = 32'h1cd712a8;
    ram_cell[   12024] = 32'h5e21101f;
    ram_cell[   12025] = 32'hda8e0dcd;
    ram_cell[   12026] = 32'hdb3e30fe;
    ram_cell[   12027] = 32'he0425389;
    ram_cell[   12028] = 32'h4c350365;
    ram_cell[   12029] = 32'habbcf020;
    ram_cell[   12030] = 32'haa106f73;
    ram_cell[   12031] = 32'h9e060908;
    ram_cell[   12032] = 32'h6657f9ff;
    ram_cell[   12033] = 32'hd64226a5;
    ram_cell[   12034] = 32'ha94d9f9c;
    ram_cell[   12035] = 32'hae8e85d1;
    ram_cell[   12036] = 32'h3601353e;
    ram_cell[   12037] = 32'h08ab6af4;
    ram_cell[   12038] = 32'h71c352a9;
    ram_cell[   12039] = 32'h66b2dd76;
    ram_cell[   12040] = 32'hf0663faa;
    ram_cell[   12041] = 32'h537b4427;
    ram_cell[   12042] = 32'he4b2a2a5;
    ram_cell[   12043] = 32'h82c392c0;
    ram_cell[   12044] = 32'h328971cd;
    ram_cell[   12045] = 32'h693af9dc;
    ram_cell[   12046] = 32'h632c19fd;
    ram_cell[   12047] = 32'h25b77b93;
    ram_cell[   12048] = 32'heb6a23d9;
    ram_cell[   12049] = 32'h2c5cbcfb;
    ram_cell[   12050] = 32'h332f994e;
    ram_cell[   12051] = 32'h1a0e208b;
    ram_cell[   12052] = 32'h24b92ee2;
    ram_cell[   12053] = 32'h271bd763;
    ram_cell[   12054] = 32'hc3254982;
    ram_cell[   12055] = 32'h58e99a04;
    ram_cell[   12056] = 32'h654fdf57;
    ram_cell[   12057] = 32'hd988dd5a;
    ram_cell[   12058] = 32'h21faa390;
    ram_cell[   12059] = 32'h3c5f5e45;
    ram_cell[   12060] = 32'h21ee4c52;
    ram_cell[   12061] = 32'h78e84271;
    ram_cell[   12062] = 32'hac53cf59;
    ram_cell[   12063] = 32'h12717c40;
    ram_cell[   12064] = 32'hcc62df96;
    ram_cell[   12065] = 32'h592884da;
    ram_cell[   12066] = 32'ha4e5ee84;
    ram_cell[   12067] = 32'h3b7456be;
    ram_cell[   12068] = 32'h03a5dedd;
    ram_cell[   12069] = 32'haf2f0a22;
    ram_cell[   12070] = 32'h22f22b5c;
    ram_cell[   12071] = 32'h777934ac;
    ram_cell[   12072] = 32'h6d634e8f;
    ram_cell[   12073] = 32'hd8138bfb;
    ram_cell[   12074] = 32'hbad706d1;
    ram_cell[   12075] = 32'h6f20fead;
    ram_cell[   12076] = 32'h334a47ed;
    ram_cell[   12077] = 32'hccb960ea;
    ram_cell[   12078] = 32'h24cafc19;
    ram_cell[   12079] = 32'he762493e;
    ram_cell[   12080] = 32'h89ce2448;
    ram_cell[   12081] = 32'h838a89ba;
    ram_cell[   12082] = 32'h4b486d97;
    ram_cell[   12083] = 32'h39a0350b;
    ram_cell[   12084] = 32'h36ee6d47;
    ram_cell[   12085] = 32'h79be71a1;
    ram_cell[   12086] = 32'h81e48c33;
    ram_cell[   12087] = 32'h7fb82a17;
    ram_cell[   12088] = 32'h3d151383;
    ram_cell[   12089] = 32'h7391ba62;
    ram_cell[   12090] = 32'h52baffb4;
    ram_cell[   12091] = 32'hc7a6e8cd;
    ram_cell[   12092] = 32'h6a367a42;
    ram_cell[   12093] = 32'hc9a55429;
    ram_cell[   12094] = 32'hc528e723;
    ram_cell[   12095] = 32'h9e566f3f;
    ram_cell[   12096] = 32'hd90a5464;
    ram_cell[   12097] = 32'h5a7b932a;
    ram_cell[   12098] = 32'h28f050e2;
    ram_cell[   12099] = 32'haab27f81;
    ram_cell[   12100] = 32'h27dc77cb;
    ram_cell[   12101] = 32'h7f3ac702;
    ram_cell[   12102] = 32'h3791b9b2;
    ram_cell[   12103] = 32'hb5b070c1;
    ram_cell[   12104] = 32'h0c2244c7;
    ram_cell[   12105] = 32'h004a490f;
    ram_cell[   12106] = 32'h6f9cd1c5;
    ram_cell[   12107] = 32'hae490b5c;
    ram_cell[   12108] = 32'hbc167e28;
    ram_cell[   12109] = 32'h177432c0;
    ram_cell[   12110] = 32'h0d48466c;
    ram_cell[   12111] = 32'hc1b155e7;
    ram_cell[   12112] = 32'h9a0031c7;
    ram_cell[   12113] = 32'hefbf34d8;
    ram_cell[   12114] = 32'h0fc51e73;
    ram_cell[   12115] = 32'h6181097e;
    ram_cell[   12116] = 32'hb031f360;
    ram_cell[   12117] = 32'h0867aae8;
    ram_cell[   12118] = 32'h1532270e;
    ram_cell[   12119] = 32'hfacbff73;
    ram_cell[   12120] = 32'ha588e9df;
    ram_cell[   12121] = 32'h6fea7468;
    ram_cell[   12122] = 32'h1ebea79b;
    ram_cell[   12123] = 32'had4a5438;
    ram_cell[   12124] = 32'h0c8dc996;
    ram_cell[   12125] = 32'h8dc39cca;
    ram_cell[   12126] = 32'hc1dc38c8;
    ram_cell[   12127] = 32'h2742f33d;
    ram_cell[   12128] = 32'hfad1a9af;
    ram_cell[   12129] = 32'h39b4d73e;
    ram_cell[   12130] = 32'h1e654b7a;
    ram_cell[   12131] = 32'h6e432eb0;
    ram_cell[   12132] = 32'he2cd302b;
    ram_cell[   12133] = 32'h522163ac;
    ram_cell[   12134] = 32'hf0ba323b;
    ram_cell[   12135] = 32'h8eb604b2;
    ram_cell[   12136] = 32'hd68bccfc;
    ram_cell[   12137] = 32'ha0484edd;
    ram_cell[   12138] = 32'h42b4dd26;
    ram_cell[   12139] = 32'heb3d3d35;
    ram_cell[   12140] = 32'h90468f2e;
    ram_cell[   12141] = 32'he9a15925;
    ram_cell[   12142] = 32'h53c36923;
    ram_cell[   12143] = 32'hbfaa0f65;
    ram_cell[   12144] = 32'hb15c6c12;
    ram_cell[   12145] = 32'ha492cb47;
    ram_cell[   12146] = 32'h810e64ca;
    ram_cell[   12147] = 32'h3c37bcb1;
    ram_cell[   12148] = 32'h046d7d52;
    ram_cell[   12149] = 32'h21cd15e8;
    ram_cell[   12150] = 32'h54dbe2ca;
    ram_cell[   12151] = 32'h793c58ff;
    ram_cell[   12152] = 32'ha558ee20;
    ram_cell[   12153] = 32'hc6bede71;
    ram_cell[   12154] = 32'h53aeaee7;
    ram_cell[   12155] = 32'h8b6c2a0e;
    ram_cell[   12156] = 32'h9ddeb007;
    ram_cell[   12157] = 32'h5fb6f274;
    ram_cell[   12158] = 32'ha42301d1;
    ram_cell[   12159] = 32'h3507bcc6;
    ram_cell[   12160] = 32'hc2406ce6;
    ram_cell[   12161] = 32'h0f30d088;
    ram_cell[   12162] = 32'hfc17907b;
    ram_cell[   12163] = 32'h55fc726d;
    ram_cell[   12164] = 32'h432f3f82;
    ram_cell[   12165] = 32'h591d9b0f;
    ram_cell[   12166] = 32'h45bca372;
    ram_cell[   12167] = 32'hba219c4c;
    ram_cell[   12168] = 32'he6a4dc34;
    ram_cell[   12169] = 32'hcfe74e50;
    ram_cell[   12170] = 32'h3bfa3753;
    ram_cell[   12171] = 32'he0b7fb35;
    ram_cell[   12172] = 32'h99899c81;
    ram_cell[   12173] = 32'h612e05b6;
    ram_cell[   12174] = 32'ha7110a5e;
    ram_cell[   12175] = 32'he6d08b14;
    ram_cell[   12176] = 32'h3db4b313;
    ram_cell[   12177] = 32'he32851a0;
    ram_cell[   12178] = 32'h52787dd0;
    ram_cell[   12179] = 32'h7a357d08;
    ram_cell[   12180] = 32'he9a483f6;
    ram_cell[   12181] = 32'h8dbcff88;
    ram_cell[   12182] = 32'h2f58bbea;
    ram_cell[   12183] = 32'h513fc978;
    ram_cell[   12184] = 32'h9a759c69;
    ram_cell[   12185] = 32'hc2533ff9;
    ram_cell[   12186] = 32'h8c1a25b6;
    ram_cell[   12187] = 32'h3ec848dc;
    ram_cell[   12188] = 32'h91f217c5;
    ram_cell[   12189] = 32'h026ffacf;
    ram_cell[   12190] = 32'h5d141620;
    ram_cell[   12191] = 32'h84b86a93;
    ram_cell[   12192] = 32'h09075b90;
    ram_cell[   12193] = 32'hc73ad319;
    ram_cell[   12194] = 32'h097b7593;
    ram_cell[   12195] = 32'h724377a4;
    ram_cell[   12196] = 32'h38ac1705;
    ram_cell[   12197] = 32'h65f15cfc;
    ram_cell[   12198] = 32'hd1d8500c;
    ram_cell[   12199] = 32'hf166cc95;
    ram_cell[   12200] = 32'he1cef150;
    ram_cell[   12201] = 32'h432a7cec;
    ram_cell[   12202] = 32'ha8fe539b;
    ram_cell[   12203] = 32'h22e2c0c3;
    ram_cell[   12204] = 32'h1fc3d710;
    ram_cell[   12205] = 32'hc28dee10;
    ram_cell[   12206] = 32'h52e1571d;
    ram_cell[   12207] = 32'hbff66604;
    ram_cell[   12208] = 32'h54732a55;
    ram_cell[   12209] = 32'h4cb9b5df;
    ram_cell[   12210] = 32'h13312499;
    ram_cell[   12211] = 32'h49ffbaf6;
    ram_cell[   12212] = 32'h1d84d3ba;
    ram_cell[   12213] = 32'ha480eabb;
    ram_cell[   12214] = 32'h89c427b4;
    ram_cell[   12215] = 32'hb174ef09;
    ram_cell[   12216] = 32'h83c168e4;
    ram_cell[   12217] = 32'h8f35c942;
    ram_cell[   12218] = 32'haafbda7f;
    ram_cell[   12219] = 32'he42c7565;
    ram_cell[   12220] = 32'hd9d0f53a;
    ram_cell[   12221] = 32'hcbcc3170;
    ram_cell[   12222] = 32'h20b4e88f;
    ram_cell[   12223] = 32'hfabdd6d8;
    ram_cell[   12224] = 32'haf2e87af;
    ram_cell[   12225] = 32'h8c2e72a8;
    ram_cell[   12226] = 32'hfa1d769a;
    ram_cell[   12227] = 32'h95d956a7;
    ram_cell[   12228] = 32'ha73075ab;
    ram_cell[   12229] = 32'hf5ffea70;
    ram_cell[   12230] = 32'hdbaf728e;
    ram_cell[   12231] = 32'h3985e6aa;
    ram_cell[   12232] = 32'h8998f9e5;
    ram_cell[   12233] = 32'hc2914249;
    ram_cell[   12234] = 32'h9fcf558c;
    ram_cell[   12235] = 32'h09ff6d7f;
    ram_cell[   12236] = 32'h021006f7;
    ram_cell[   12237] = 32'hded29fa2;
    ram_cell[   12238] = 32'h7966590f;
    ram_cell[   12239] = 32'hf37ed7dc;
    ram_cell[   12240] = 32'hf18aa56d;
    ram_cell[   12241] = 32'h6a0387f0;
    ram_cell[   12242] = 32'h47f02039;
    ram_cell[   12243] = 32'h6eb4bbc1;
    ram_cell[   12244] = 32'h7015709a;
    ram_cell[   12245] = 32'h46fe6be4;
    ram_cell[   12246] = 32'h17f6e8f0;
    ram_cell[   12247] = 32'h080cf2a2;
    ram_cell[   12248] = 32'h3d6f745e;
    ram_cell[   12249] = 32'h46c19985;
    ram_cell[   12250] = 32'h553251fa;
    ram_cell[   12251] = 32'h4f3ed83d;
    ram_cell[   12252] = 32'h4996ca8c;
    ram_cell[   12253] = 32'h68e07854;
    ram_cell[   12254] = 32'h6d9d1ad4;
    ram_cell[   12255] = 32'h6b97103d;
    ram_cell[   12256] = 32'h4ea5411f;
    ram_cell[   12257] = 32'h7b5189d0;
    ram_cell[   12258] = 32'h7d0fdfa2;
    ram_cell[   12259] = 32'h492d0fa2;
    ram_cell[   12260] = 32'hfdd781ec;
    ram_cell[   12261] = 32'h89667eae;
    ram_cell[   12262] = 32'h69cea9e0;
    ram_cell[   12263] = 32'h52498724;
    ram_cell[   12264] = 32'h7d42b780;
    ram_cell[   12265] = 32'he3e9b7b6;
    ram_cell[   12266] = 32'hfd712b66;
    ram_cell[   12267] = 32'h52a814f7;
    ram_cell[   12268] = 32'h5e110ad9;
    ram_cell[   12269] = 32'h8c25d7da;
    ram_cell[   12270] = 32'hc22c50b8;
    ram_cell[   12271] = 32'h899ea0de;
    ram_cell[   12272] = 32'hfa23a314;
    ram_cell[   12273] = 32'hbacc6699;
    ram_cell[   12274] = 32'hebf51739;
    ram_cell[   12275] = 32'h39ea4186;
    ram_cell[   12276] = 32'hcbc809d3;
    ram_cell[   12277] = 32'hffc25347;
    ram_cell[   12278] = 32'hac5dab36;
    ram_cell[   12279] = 32'he055a1f0;
    ram_cell[   12280] = 32'hb21d76c8;
    ram_cell[   12281] = 32'h31ede7bc;
    ram_cell[   12282] = 32'h6bb05b00;
    ram_cell[   12283] = 32'hfda54c90;
    ram_cell[   12284] = 32'h75a2bbbb;
    ram_cell[   12285] = 32'h89a0240d;
    ram_cell[   12286] = 32'h5ec613e7;
    ram_cell[   12287] = 32'hbf222be9;
end

endmodule

