
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'haadda71b;
    ram_cell[       1] = 32'h0;  // 32'h58816d4c;
    ram_cell[       2] = 32'h0;  // 32'h6329fa82;
    ram_cell[       3] = 32'h0;  // 32'h7dca74f6;
    ram_cell[       4] = 32'h0;  // 32'hd955bc4b;
    ram_cell[       5] = 32'h0;  // 32'hc24faae6;
    ram_cell[       6] = 32'h0;  // 32'he600d5e9;
    ram_cell[       7] = 32'h0;  // 32'h2576a220;
    ram_cell[       8] = 32'h0;  // 32'h8b532999;
    ram_cell[       9] = 32'h0;  // 32'hb2e49081;
    ram_cell[      10] = 32'h0;  // 32'hdcdf90c6;
    ram_cell[      11] = 32'h0;  // 32'h4f20cc82;
    ram_cell[      12] = 32'h0;  // 32'h6313eb6f;
    ram_cell[      13] = 32'h0;  // 32'h9dc44d2b;
    ram_cell[      14] = 32'h0;  // 32'h7f3b240c;
    ram_cell[      15] = 32'h0;  // 32'h2411b667;
    ram_cell[      16] = 32'h0;  // 32'hade56d5e;
    ram_cell[      17] = 32'h0;  // 32'ha7fcc157;
    ram_cell[      18] = 32'h0;  // 32'hc7107940;
    ram_cell[      19] = 32'h0;  // 32'h931ff246;
    ram_cell[      20] = 32'h0;  // 32'h6bc0cd6b;
    ram_cell[      21] = 32'h0;  // 32'h4ac6ea19;
    ram_cell[      22] = 32'h0;  // 32'hb0e3cc41;
    ram_cell[      23] = 32'h0;  // 32'h2f395761;
    ram_cell[      24] = 32'h0;  // 32'ha7287ef0;
    ram_cell[      25] = 32'h0;  // 32'h66d2c613;
    ram_cell[      26] = 32'h0;  // 32'h5b6875c9;
    ram_cell[      27] = 32'h0;  // 32'hb7cd0314;
    ram_cell[      28] = 32'h0;  // 32'hfc81dd01;
    ram_cell[      29] = 32'h0;  // 32'h582f737f;
    ram_cell[      30] = 32'h0;  // 32'h8ee296f7;
    ram_cell[      31] = 32'h0;  // 32'h052833de;
    ram_cell[      32] = 32'h0;  // 32'hb1824a10;
    ram_cell[      33] = 32'h0;  // 32'hd61ae49c;
    ram_cell[      34] = 32'h0;  // 32'hd1687c89;
    ram_cell[      35] = 32'h0;  // 32'h302038d7;
    ram_cell[      36] = 32'h0;  // 32'hdad67321;
    ram_cell[      37] = 32'h0;  // 32'he1f112ca;
    ram_cell[      38] = 32'h0;  // 32'hd24afd98;
    ram_cell[      39] = 32'h0;  // 32'hdd8d72e3;
    ram_cell[      40] = 32'h0;  // 32'h81dc8f4e;
    ram_cell[      41] = 32'h0;  // 32'hdb6109cc;
    ram_cell[      42] = 32'h0;  // 32'h882fffcd;
    ram_cell[      43] = 32'h0;  // 32'h645e4e50;
    ram_cell[      44] = 32'h0;  // 32'h067b0974;
    ram_cell[      45] = 32'h0;  // 32'ha6a10d11;
    ram_cell[      46] = 32'h0;  // 32'h8a4c20e6;
    ram_cell[      47] = 32'h0;  // 32'he50ba0cc;
    ram_cell[      48] = 32'h0;  // 32'hdcbb2398;
    ram_cell[      49] = 32'h0;  // 32'h5ba7e78f;
    ram_cell[      50] = 32'h0;  // 32'h5abe1f0f;
    ram_cell[      51] = 32'h0;  // 32'ha34a62dc;
    ram_cell[      52] = 32'h0;  // 32'h46369067;
    ram_cell[      53] = 32'h0;  // 32'h2e089877;
    ram_cell[      54] = 32'h0;  // 32'hcb74adbb;
    ram_cell[      55] = 32'h0;  // 32'he1fac2d6;
    ram_cell[      56] = 32'h0;  // 32'h93e98cbc;
    ram_cell[      57] = 32'h0;  // 32'h68a1e28a;
    ram_cell[      58] = 32'h0;  // 32'hce956098;
    ram_cell[      59] = 32'h0;  // 32'hee51a401;
    ram_cell[      60] = 32'h0;  // 32'h569cc656;
    ram_cell[      61] = 32'h0;  // 32'h158db5a7;
    ram_cell[      62] = 32'h0;  // 32'h9394d376;
    ram_cell[      63] = 32'h0;  // 32'hda84224d;
    ram_cell[      64] = 32'h0;  // 32'hea0247ec;
    ram_cell[      65] = 32'h0;  // 32'h9db1430c;
    ram_cell[      66] = 32'h0;  // 32'h6fff0e60;
    ram_cell[      67] = 32'h0;  // 32'h29a41f6d;
    ram_cell[      68] = 32'h0;  // 32'hc0532987;
    ram_cell[      69] = 32'h0;  // 32'h6cfb672e;
    ram_cell[      70] = 32'h0;  // 32'h5712e738;
    ram_cell[      71] = 32'h0;  // 32'h0cfe90c9;
    ram_cell[      72] = 32'h0;  // 32'h54aa032e;
    ram_cell[      73] = 32'h0;  // 32'hdef7aa07;
    ram_cell[      74] = 32'h0;  // 32'hfbe38893;
    ram_cell[      75] = 32'h0;  // 32'h4f6a70d8;
    ram_cell[      76] = 32'h0;  // 32'hbb780e1a;
    ram_cell[      77] = 32'h0;  // 32'he8eea142;
    ram_cell[      78] = 32'h0;  // 32'h4bce3f0b;
    ram_cell[      79] = 32'h0;  // 32'hc351acbc;
    ram_cell[      80] = 32'h0;  // 32'h67a8957d;
    ram_cell[      81] = 32'h0;  // 32'h1339e146;
    ram_cell[      82] = 32'h0;  // 32'h19597c78;
    ram_cell[      83] = 32'h0;  // 32'h27bc3b09;
    ram_cell[      84] = 32'h0;  // 32'h5d16e553;
    ram_cell[      85] = 32'h0;  // 32'h5ef074b0;
    ram_cell[      86] = 32'h0;  // 32'hf7d701e3;
    ram_cell[      87] = 32'h0;  // 32'h29355cd0;
    ram_cell[      88] = 32'h0;  // 32'hc77ca219;
    ram_cell[      89] = 32'h0;  // 32'h01ccf07d;
    ram_cell[      90] = 32'h0;  // 32'ha645af9c;
    ram_cell[      91] = 32'h0;  // 32'hd2853765;
    ram_cell[      92] = 32'h0;  // 32'h4e0079bb;
    ram_cell[      93] = 32'h0;  // 32'he1e1e970;
    ram_cell[      94] = 32'h0;  // 32'h3ab03edf;
    ram_cell[      95] = 32'h0;  // 32'h728337c1;
    ram_cell[      96] = 32'h0;  // 32'h778195b3;
    ram_cell[      97] = 32'h0;  // 32'hd065436b;
    ram_cell[      98] = 32'h0;  // 32'hb41f06d7;
    ram_cell[      99] = 32'h0;  // 32'h41bea69d;
    ram_cell[     100] = 32'h0;  // 32'h6d398c65;
    ram_cell[     101] = 32'h0;  // 32'h11739b9d;
    ram_cell[     102] = 32'h0;  // 32'h7fde18f1;
    ram_cell[     103] = 32'h0;  // 32'hc845239d;
    ram_cell[     104] = 32'h0;  // 32'h35f1d386;
    ram_cell[     105] = 32'h0;  // 32'hb3ab288b;
    ram_cell[     106] = 32'h0;  // 32'h767ae90e;
    ram_cell[     107] = 32'h0;  // 32'h953ff056;
    ram_cell[     108] = 32'h0;  // 32'hc2f931cc;
    ram_cell[     109] = 32'h0;  // 32'h2a9eb3bc;
    ram_cell[     110] = 32'h0;  // 32'h562d3510;
    ram_cell[     111] = 32'h0;  // 32'h23c2ec88;
    ram_cell[     112] = 32'h0;  // 32'hbcf7f64a;
    ram_cell[     113] = 32'h0;  // 32'h9b39bc0a;
    ram_cell[     114] = 32'h0;  // 32'h8940fe0b;
    ram_cell[     115] = 32'h0;  // 32'hbc67fe80;
    ram_cell[     116] = 32'h0;  // 32'hcb84959a;
    ram_cell[     117] = 32'h0;  // 32'hcc0b7e9f;
    ram_cell[     118] = 32'h0;  // 32'hfa757359;
    ram_cell[     119] = 32'h0;  // 32'hee5eec62;
    ram_cell[     120] = 32'h0;  // 32'haa864721;
    ram_cell[     121] = 32'h0;  // 32'h9c44a4d0;
    ram_cell[     122] = 32'h0;  // 32'hde384662;
    ram_cell[     123] = 32'h0;  // 32'h67bb8b09;
    ram_cell[     124] = 32'h0;  // 32'h2d40b7fc;
    ram_cell[     125] = 32'h0;  // 32'hc8802e8b;
    ram_cell[     126] = 32'h0;  // 32'hd88213b4;
    ram_cell[     127] = 32'h0;  // 32'h5c627fc8;
    ram_cell[     128] = 32'h0;  // 32'h4c745dfb;
    ram_cell[     129] = 32'h0;  // 32'h8fd82c40;
    ram_cell[     130] = 32'h0;  // 32'h30a4d782;
    ram_cell[     131] = 32'h0;  // 32'h2c28c6cc;
    ram_cell[     132] = 32'h0;  // 32'h5aba1dd7;
    ram_cell[     133] = 32'h0;  // 32'h85ac86d7;
    ram_cell[     134] = 32'h0;  // 32'hc1de3dbf;
    ram_cell[     135] = 32'h0;  // 32'h7cedab31;
    ram_cell[     136] = 32'h0;  // 32'hec59892f;
    ram_cell[     137] = 32'h0;  // 32'h730e7aed;
    ram_cell[     138] = 32'h0;  // 32'h274812e2;
    ram_cell[     139] = 32'h0;  // 32'hb8c643cf;
    ram_cell[     140] = 32'h0;  // 32'haa27796b;
    ram_cell[     141] = 32'h0;  // 32'hb3ec97b9;
    ram_cell[     142] = 32'h0;  // 32'h711552f4;
    ram_cell[     143] = 32'h0;  // 32'h1f8c8976;
    ram_cell[     144] = 32'h0;  // 32'h5cbc698f;
    ram_cell[     145] = 32'h0;  // 32'h4f892ceb;
    ram_cell[     146] = 32'h0;  // 32'h1d43c2d3;
    ram_cell[     147] = 32'h0;  // 32'h0bce3967;
    ram_cell[     148] = 32'h0;  // 32'h2bb79a21;
    ram_cell[     149] = 32'h0;  // 32'he2039fe2;
    ram_cell[     150] = 32'h0;  // 32'h479b368a;
    ram_cell[     151] = 32'h0;  // 32'h7b8cb974;
    ram_cell[     152] = 32'h0;  // 32'hcd7c6872;
    ram_cell[     153] = 32'h0;  // 32'hf2530c21;
    ram_cell[     154] = 32'h0;  // 32'hfa551275;
    ram_cell[     155] = 32'h0;  // 32'hfeefab37;
    ram_cell[     156] = 32'h0;  // 32'h924c0fc3;
    ram_cell[     157] = 32'h0;  // 32'ha41b6f2c;
    ram_cell[     158] = 32'h0;  // 32'hd117b728;
    ram_cell[     159] = 32'h0;  // 32'h0b7ff83d;
    ram_cell[     160] = 32'h0;  // 32'h58b25b2c;
    ram_cell[     161] = 32'h0;  // 32'h5781cee3;
    ram_cell[     162] = 32'h0;  // 32'hff8aea80;
    ram_cell[     163] = 32'h0;  // 32'hf38508ab;
    ram_cell[     164] = 32'h0;  // 32'hea9a192b;
    ram_cell[     165] = 32'h0;  // 32'hb3b89309;
    ram_cell[     166] = 32'h0;  // 32'h5890d49b;
    ram_cell[     167] = 32'h0;  // 32'h93ded848;
    ram_cell[     168] = 32'h0;  // 32'h74473333;
    ram_cell[     169] = 32'h0;  // 32'hd45d9fc3;
    ram_cell[     170] = 32'h0;  // 32'h6f331b5c;
    ram_cell[     171] = 32'h0;  // 32'hb76f8588;
    ram_cell[     172] = 32'h0;  // 32'he165314d;
    ram_cell[     173] = 32'h0;  // 32'h5cd26619;
    ram_cell[     174] = 32'h0;  // 32'hdb0b2049;
    ram_cell[     175] = 32'h0;  // 32'hcdb4e62e;
    ram_cell[     176] = 32'h0;  // 32'hd1fbf813;
    ram_cell[     177] = 32'h0;  // 32'h16ef932b;
    ram_cell[     178] = 32'h0;  // 32'h99e3e40c;
    ram_cell[     179] = 32'h0;  // 32'h969226a8;
    ram_cell[     180] = 32'h0;  // 32'h87f57ffe;
    ram_cell[     181] = 32'h0;  // 32'h0bc050e2;
    ram_cell[     182] = 32'h0;  // 32'h9cb31219;
    ram_cell[     183] = 32'h0;  // 32'h4fec2027;
    ram_cell[     184] = 32'h0;  // 32'h069407fd;
    ram_cell[     185] = 32'h0;  // 32'ha12bed4e;
    ram_cell[     186] = 32'h0;  // 32'h5bb62e7a;
    ram_cell[     187] = 32'h0;  // 32'h94b3cf9c;
    ram_cell[     188] = 32'h0;  // 32'hd6a3bdd0;
    ram_cell[     189] = 32'h0;  // 32'hce96c4a4;
    ram_cell[     190] = 32'h0;  // 32'h30bb85b2;
    ram_cell[     191] = 32'h0;  // 32'hf0603c1d;
    ram_cell[     192] = 32'h0;  // 32'h9c9e88cc;
    ram_cell[     193] = 32'h0;  // 32'h4f9d661b;
    ram_cell[     194] = 32'h0;  // 32'hb951e28e;
    ram_cell[     195] = 32'h0;  // 32'he2e60ae3;
    ram_cell[     196] = 32'h0;  // 32'hc62a1f68;
    ram_cell[     197] = 32'h0;  // 32'h828bb0f6;
    ram_cell[     198] = 32'h0;  // 32'h9308523b;
    ram_cell[     199] = 32'h0;  // 32'h18000278;
    ram_cell[     200] = 32'h0;  // 32'h22adc8b3;
    ram_cell[     201] = 32'h0;  // 32'h4d0789c5;
    ram_cell[     202] = 32'h0;  // 32'h8e5f2055;
    ram_cell[     203] = 32'h0;  // 32'h74faf71f;
    ram_cell[     204] = 32'h0;  // 32'h6a372735;
    ram_cell[     205] = 32'h0;  // 32'h89ced6a9;
    ram_cell[     206] = 32'h0;  // 32'h12b58bdd;
    ram_cell[     207] = 32'h0;  // 32'h6014b01a;
    ram_cell[     208] = 32'h0;  // 32'h6d1abe8b;
    ram_cell[     209] = 32'h0;  // 32'h425dc0e2;
    ram_cell[     210] = 32'h0;  // 32'h16c476ca;
    ram_cell[     211] = 32'h0;  // 32'h4648a112;
    ram_cell[     212] = 32'h0;  // 32'h93e66deb;
    ram_cell[     213] = 32'h0;  // 32'h7f9f38a4;
    ram_cell[     214] = 32'h0;  // 32'h6cc601c8;
    ram_cell[     215] = 32'h0;  // 32'hfeff6a26;
    ram_cell[     216] = 32'h0;  // 32'hd29a0d75;
    ram_cell[     217] = 32'h0;  // 32'h6d412127;
    ram_cell[     218] = 32'h0;  // 32'h1385a21b;
    ram_cell[     219] = 32'h0;  // 32'hc8384031;
    ram_cell[     220] = 32'h0;  // 32'hd657c24a;
    ram_cell[     221] = 32'h0;  // 32'h51bae8fe;
    ram_cell[     222] = 32'h0;  // 32'h1c3daa5b;
    ram_cell[     223] = 32'h0;  // 32'h21115056;
    ram_cell[     224] = 32'h0;  // 32'h32151533;
    ram_cell[     225] = 32'h0;  // 32'haa9fdf4b;
    ram_cell[     226] = 32'h0;  // 32'hfdd0bf59;
    ram_cell[     227] = 32'h0;  // 32'h8051c9be;
    ram_cell[     228] = 32'h0;  // 32'hb1aef71b;
    ram_cell[     229] = 32'h0;  // 32'h806470d1;
    ram_cell[     230] = 32'h0;  // 32'h87c569df;
    ram_cell[     231] = 32'h0;  // 32'haaf89c02;
    ram_cell[     232] = 32'h0;  // 32'h3c2c88f5;
    ram_cell[     233] = 32'h0;  // 32'h70302596;
    ram_cell[     234] = 32'h0;  // 32'h870db486;
    ram_cell[     235] = 32'h0;  // 32'h783ec424;
    ram_cell[     236] = 32'h0;  // 32'h113c5ffc;
    ram_cell[     237] = 32'h0;  // 32'h138d4e6d;
    ram_cell[     238] = 32'h0;  // 32'h1669dd52;
    ram_cell[     239] = 32'h0;  // 32'h72e58d25;
    ram_cell[     240] = 32'h0;  // 32'h831a3f35;
    ram_cell[     241] = 32'h0;  // 32'hc22155f5;
    ram_cell[     242] = 32'h0;  // 32'h931c8ccf;
    ram_cell[     243] = 32'h0;  // 32'ha238be4a;
    ram_cell[     244] = 32'h0;  // 32'h16deb447;
    ram_cell[     245] = 32'h0;  // 32'h9f6b4d9c;
    ram_cell[     246] = 32'h0;  // 32'h71facdf9;
    ram_cell[     247] = 32'h0;  // 32'h62487730;
    ram_cell[     248] = 32'h0;  // 32'hbd4b9806;
    ram_cell[     249] = 32'h0;  // 32'hd0e0bc5d;
    ram_cell[     250] = 32'h0;  // 32'h3de566b5;
    ram_cell[     251] = 32'h0;  // 32'hd220a3d7;
    ram_cell[     252] = 32'h0;  // 32'h5df9afb8;
    ram_cell[     253] = 32'h0;  // 32'hdeeadaf6;
    ram_cell[     254] = 32'h0;  // 32'ha8eb08f7;
    ram_cell[     255] = 32'h0;  // 32'h0ddb1d28;
    // src matrix A
    ram_cell[     256] = 32'hff3d7e65;
    ram_cell[     257] = 32'hbf26fab4;
    ram_cell[     258] = 32'h29bfde49;
    ram_cell[     259] = 32'h8f2e697e;
    ram_cell[     260] = 32'h49c07c13;
    ram_cell[     261] = 32'hb276b4c3;
    ram_cell[     262] = 32'h06396047;
    ram_cell[     263] = 32'h13db785e;
    ram_cell[     264] = 32'h66896259;
    ram_cell[     265] = 32'h03d00a54;
    ram_cell[     266] = 32'hfa1e480b;
    ram_cell[     267] = 32'h496068e8;
    ram_cell[     268] = 32'h497181ba;
    ram_cell[     269] = 32'he2571558;
    ram_cell[     270] = 32'ha7a6c678;
    ram_cell[     271] = 32'h9582d8ee;
    ram_cell[     272] = 32'h151e2472;
    ram_cell[     273] = 32'h5934934c;
    ram_cell[     274] = 32'h8a34cb4c;
    ram_cell[     275] = 32'hbfbb6de4;
    ram_cell[     276] = 32'h3a7dc054;
    ram_cell[     277] = 32'h299f1952;
    ram_cell[     278] = 32'ha485b85c;
    ram_cell[     279] = 32'h854259dc;
    ram_cell[     280] = 32'h5d2269a7;
    ram_cell[     281] = 32'h143e6a6a;
    ram_cell[     282] = 32'h25c46dae;
    ram_cell[     283] = 32'h732d4954;
    ram_cell[     284] = 32'h9dda8bc3;
    ram_cell[     285] = 32'h78681565;
    ram_cell[     286] = 32'h37678894;
    ram_cell[     287] = 32'h26138490;
    ram_cell[     288] = 32'h8521876e;
    ram_cell[     289] = 32'he631d562;
    ram_cell[     290] = 32'hf4b42df9;
    ram_cell[     291] = 32'hd44357a1;
    ram_cell[     292] = 32'h568b7acc;
    ram_cell[     293] = 32'h1803e513;
    ram_cell[     294] = 32'h4eaa9898;
    ram_cell[     295] = 32'h4b4e360e;
    ram_cell[     296] = 32'he98b4679;
    ram_cell[     297] = 32'h85339541;
    ram_cell[     298] = 32'h54a4535e;
    ram_cell[     299] = 32'hd715f1c3;
    ram_cell[     300] = 32'hd6c5a65e;
    ram_cell[     301] = 32'h18798a31;
    ram_cell[     302] = 32'hef9120f8;
    ram_cell[     303] = 32'ha0824b8c;
    ram_cell[     304] = 32'h62c03744;
    ram_cell[     305] = 32'h4ef7d666;
    ram_cell[     306] = 32'haaa57b7e;
    ram_cell[     307] = 32'h9775b764;
    ram_cell[     308] = 32'ha16284eb;
    ram_cell[     309] = 32'h6f586fd6;
    ram_cell[     310] = 32'h3a5bed2d;
    ram_cell[     311] = 32'h5003c209;
    ram_cell[     312] = 32'h3aa72054;
    ram_cell[     313] = 32'h8427afe8;
    ram_cell[     314] = 32'h30692cd7;
    ram_cell[     315] = 32'h16595416;
    ram_cell[     316] = 32'ha74eba4c;
    ram_cell[     317] = 32'h971bfe53;
    ram_cell[     318] = 32'hbdde1820;
    ram_cell[     319] = 32'h13f3aa31;
    ram_cell[     320] = 32'h7125426f;
    ram_cell[     321] = 32'he91974ef;
    ram_cell[     322] = 32'h26735af5;
    ram_cell[     323] = 32'hb4702c52;
    ram_cell[     324] = 32'hb6d37256;
    ram_cell[     325] = 32'he5eaf8cf;
    ram_cell[     326] = 32'h12e1d79b;
    ram_cell[     327] = 32'h6f540bb9;
    ram_cell[     328] = 32'hf3fb3286;
    ram_cell[     329] = 32'h248c06e5;
    ram_cell[     330] = 32'hb1c1543e;
    ram_cell[     331] = 32'h1d1c21f1;
    ram_cell[     332] = 32'h40fd2f25;
    ram_cell[     333] = 32'h116ce019;
    ram_cell[     334] = 32'h0b00f0c6;
    ram_cell[     335] = 32'h06c63ec4;
    ram_cell[     336] = 32'h54867e10;
    ram_cell[     337] = 32'h3b94bbbc;
    ram_cell[     338] = 32'h72d7fc40;
    ram_cell[     339] = 32'h19c47bb2;
    ram_cell[     340] = 32'h8c187f43;
    ram_cell[     341] = 32'h61405af7;
    ram_cell[     342] = 32'h97e79b98;
    ram_cell[     343] = 32'ha0afaeee;
    ram_cell[     344] = 32'hc268136e;
    ram_cell[     345] = 32'h565db200;
    ram_cell[     346] = 32'hed1f527e;
    ram_cell[     347] = 32'h1d2234ae;
    ram_cell[     348] = 32'h75f8d21e;
    ram_cell[     349] = 32'h3620bffb;
    ram_cell[     350] = 32'h08c3fc75;
    ram_cell[     351] = 32'hd3cf662a;
    ram_cell[     352] = 32'h2cdbc53f;
    ram_cell[     353] = 32'h347b11df;
    ram_cell[     354] = 32'h296e9c32;
    ram_cell[     355] = 32'h95bd5c58;
    ram_cell[     356] = 32'had680f17;
    ram_cell[     357] = 32'hb0a3f694;
    ram_cell[     358] = 32'h7f361621;
    ram_cell[     359] = 32'hbc191815;
    ram_cell[     360] = 32'h5f11eba8;
    ram_cell[     361] = 32'h722fe373;
    ram_cell[     362] = 32'h44fbd831;
    ram_cell[     363] = 32'h801930ec;
    ram_cell[     364] = 32'hc01a35f6;
    ram_cell[     365] = 32'h7d7a55b0;
    ram_cell[     366] = 32'hf4c8922b;
    ram_cell[     367] = 32'hc6ecd880;
    ram_cell[     368] = 32'he5493fc0;
    ram_cell[     369] = 32'h2bb2b8cb;
    ram_cell[     370] = 32'hf5719085;
    ram_cell[     371] = 32'h5531d404;
    ram_cell[     372] = 32'h83bf9192;
    ram_cell[     373] = 32'h126a3e04;
    ram_cell[     374] = 32'hd2fb3250;
    ram_cell[     375] = 32'h8d906dd8;
    ram_cell[     376] = 32'h44c7ce20;
    ram_cell[     377] = 32'h6389026a;
    ram_cell[     378] = 32'h493f7bf9;
    ram_cell[     379] = 32'hda6a8587;
    ram_cell[     380] = 32'h448ca41f;
    ram_cell[     381] = 32'h7ee2c396;
    ram_cell[     382] = 32'h1f531218;
    ram_cell[     383] = 32'h48ae1eba;
    ram_cell[     384] = 32'h11d63eb7;
    ram_cell[     385] = 32'hb994c2b5;
    ram_cell[     386] = 32'hcc20d39a;
    ram_cell[     387] = 32'hb702e305;
    ram_cell[     388] = 32'hbc92b81c;
    ram_cell[     389] = 32'h67051331;
    ram_cell[     390] = 32'hde0c80d8;
    ram_cell[     391] = 32'h22e26658;
    ram_cell[     392] = 32'hb2ee3dc4;
    ram_cell[     393] = 32'h1786ef3f;
    ram_cell[     394] = 32'h27d0f97a;
    ram_cell[     395] = 32'hbbe0884a;
    ram_cell[     396] = 32'ha8a3c23d;
    ram_cell[     397] = 32'h709ca2e5;
    ram_cell[     398] = 32'h080dbee5;
    ram_cell[     399] = 32'h96926a51;
    ram_cell[     400] = 32'h127a40dc;
    ram_cell[     401] = 32'h4717dda6;
    ram_cell[     402] = 32'h06e8f47e;
    ram_cell[     403] = 32'h957a7c2e;
    ram_cell[     404] = 32'h09686a35;
    ram_cell[     405] = 32'h30f5d77c;
    ram_cell[     406] = 32'hac11838d;
    ram_cell[     407] = 32'h90e5623c;
    ram_cell[     408] = 32'he18953d3;
    ram_cell[     409] = 32'h2bf85c89;
    ram_cell[     410] = 32'h0887ea28;
    ram_cell[     411] = 32'h849e99f2;
    ram_cell[     412] = 32'hd9188d9c;
    ram_cell[     413] = 32'hea4d670a;
    ram_cell[     414] = 32'h0d6b78a9;
    ram_cell[     415] = 32'h7f69db98;
    ram_cell[     416] = 32'he2df2aef;
    ram_cell[     417] = 32'h84502ff4;
    ram_cell[     418] = 32'ha82870ff;
    ram_cell[     419] = 32'hda84fa15;
    ram_cell[     420] = 32'hc7ea647e;
    ram_cell[     421] = 32'h96fb5c1f;
    ram_cell[     422] = 32'h8b9acffe;
    ram_cell[     423] = 32'ha29c5af1;
    ram_cell[     424] = 32'h3b2b6d8e;
    ram_cell[     425] = 32'h72d3319e;
    ram_cell[     426] = 32'hd0e0362b;
    ram_cell[     427] = 32'h6698d00f;
    ram_cell[     428] = 32'he80bc4c7;
    ram_cell[     429] = 32'he02b9ab0;
    ram_cell[     430] = 32'h38e74726;
    ram_cell[     431] = 32'h4e16fd5e;
    ram_cell[     432] = 32'h04db1901;
    ram_cell[     433] = 32'hafde6d43;
    ram_cell[     434] = 32'h29bde598;
    ram_cell[     435] = 32'h20ac70b9;
    ram_cell[     436] = 32'h3974c88d;
    ram_cell[     437] = 32'h08cbccf6;
    ram_cell[     438] = 32'h2c9aa7e6;
    ram_cell[     439] = 32'ha496200e;
    ram_cell[     440] = 32'had89322c;
    ram_cell[     441] = 32'hd88643ab;
    ram_cell[     442] = 32'hba957bc9;
    ram_cell[     443] = 32'he845b1df;
    ram_cell[     444] = 32'h00cbdc24;
    ram_cell[     445] = 32'h0b883df7;
    ram_cell[     446] = 32'hd4739e94;
    ram_cell[     447] = 32'hde3ffe86;
    ram_cell[     448] = 32'hf5a17266;
    ram_cell[     449] = 32'h200371af;
    ram_cell[     450] = 32'h31ef3f65;
    ram_cell[     451] = 32'h06249b01;
    ram_cell[     452] = 32'h5b58fc67;
    ram_cell[     453] = 32'h91d658cf;
    ram_cell[     454] = 32'hcc971e14;
    ram_cell[     455] = 32'h6fd0d153;
    ram_cell[     456] = 32'hb0517f01;
    ram_cell[     457] = 32'h24c20a4e;
    ram_cell[     458] = 32'h67950a98;
    ram_cell[     459] = 32'h323137a7;
    ram_cell[     460] = 32'h83dd6f6e;
    ram_cell[     461] = 32'ha540f22b;
    ram_cell[     462] = 32'h2851cd15;
    ram_cell[     463] = 32'h6618bc36;
    ram_cell[     464] = 32'h05d490ea;
    ram_cell[     465] = 32'h081ff9ea;
    ram_cell[     466] = 32'hf4459cb6;
    ram_cell[     467] = 32'hfc4219cc;
    ram_cell[     468] = 32'h3ee3d1a1;
    ram_cell[     469] = 32'hfe0487d4;
    ram_cell[     470] = 32'h3ca30f5f;
    ram_cell[     471] = 32'h57bc3bd1;
    ram_cell[     472] = 32'h6a462459;
    ram_cell[     473] = 32'he45cc5ff;
    ram_cell[     474] = 32'h8d395ea2;
    ram_cell[     475] = 32'h7c7a7367;
    ram_cell[     476] = 32'h434831c5;
    ram_cell[     477] = 32'h569d2273;
    ram_cell[     478] = 32'h59d6e2e4;
    ram_cell[     479] = 32'ha769d7a6;
    ram_cell[     480] = 32'h553d7c41;
    ram_cell[     481] = 32'h64e2cb88;
    ram_cell[     482] = 32'h9de0cf7b;
    ram_cell[     483] = 32'haae784df;
    ram_cell[     484] = 32'h7c7ae0e6;
    ram_cell[     485] = 32'hd6c6919c;
    ram_cell[     486] = 32'hcee3cf4d;
    ram_cell[     487] = 32'he70440cc;
    ram_cell[     488] = 32'h82e1e8db;
    ram_cell[     489] = 32'hb09a7625;
    ram_cell[     490] = 32'hd75fd212;
    ram_cell[     491] = 32'he0732221;
    ram_cell[     492] = 32'hc83a2fd4;
    ram_cell[     493] = 32'h10d0d27a;
    ram_cell[     494] = 32'hf974bbd9;
    ram_cell[     495] = 32'h1e91a7a8;
    ram_cell[     496] = 32'h4f030717;
    ram_cell[     497] = 32'hba19f5bf;
    ram_cell[     498] = 32'h0203cdc0;
    ram_cell[     499] = 32'h0475ee7d;
    ram_cell[     500] = 32'he6abc06d;
    ram_cell[     501] = 32'he71f1564;
    ram_cell[     502] = 32'hf56acb54;
    ram_cell[     503] = 32'h5a8748fc;
    ram_cell[     504] = 32'hd6cc2e91;
    ram_cell[     505] = 32'hda847256;
    ram_cell[     506] = 32'h0eee9043;
    ram_cell[     507] = 32'hba612125;
    ram_cell[     508] = 32'h75882673;
    ram_cell[     509] = 32'hbabcb664;
    ram_cell[     510] = 32'h2c142468;
    ram_cell[     511] = 32'hbd6dcbae;
    // src matrix B
    ram_cell[     512] = 32'h4f57e8b7;
    ram_cell[     513] = 32'h9e897f6f;
    ram_cell[     514] = 32'h9b480b0c;
    ram_cell[     515] = 32'hdb3aa5c7;
    ram_cell[     516] = 32'h97ce21ba;
    ram_cell[     517] = 32'h6a63afc9;
    ram_cell[     518] = 32'h491b34b6;
    ram_cell[     519] = 32'he65073bd;
    ram_cell[     520] = 32'h36d9c3f9;
    ram_cell[     521] = 32'h9152a798;
    ram_cell[     522] = 32'h10ff40c7;
    ram_cell[     523] = 32'h813a09dc;
    ram_cell[     524] = 32'hbeeafea1;
    ram_cell[     525] = 32'h01982fa2;
    ram_cell[     526] = 32'hbf9a8ded;
    ram_cell[     527] = 32'h95a0d160;
    ram_cell[     528] = 32'h18416ad2;
    ram_cell[     529] = 32'hd1160975;
    ram_cell[     530] = 32'h04d68ef6;
    ram_cell[     531] = 32'h44c016f7;
    ram_cell[     532] = 32'h8914531b;
    ram_cell[     533] = 32'h7e044d36;
    ram_cell[     534] = 32'h025d06a7;
    ram_cell[     535] = 32'hf006ea48;
    ram_cell[     536] = 32'hfc5483c4;
    ram_cell[     537] = 32'hac490aed;
    ram_cell[     538] = 32'hcbb39fe3;
    ram_cell[     539] = 32'h95cf9282;
    ram_cell[     540] = 32'h1216b479;
    ram_cell[     541] = 32'h1ae3f797;
    ram_cell[     542] = 32'h7f7df912;
    ram_cell[     543] = 32'h8895bc39;
    ram_cell[     544] = 32'h102c7c89;
    ram_cell[     545] = 32'h7920bfaf;
    ram_cell[     546] = 32'h02832752;
    ram_cell[     547] = 32'h2fa129cc;
    ram_cell[     548] = 32'h707d7b66;
    ram_cell[     549] = 32'h11158ff3;
    ram_cell[     550] = 32'hcb59e8d1;
    ram_cell[     551] = 32'hb86b31c9;
    ram_cell[     552] = 32'h44e6e832;
    ram_cell[     553] = 32'h2ba44d14;
    ram_cell[     554] = 32'h003905b0;
    ram_cell[     555] = 32'ha6d6a9aa;
    ram_cell[     556] = 32'h03d1bf57;
    ram_cell[     557] = 32'hdbab9ffa;
    ram_cell[     558] = 32'h0962b340;
    ram_cell[     559] = 32'hdf242681;
    ram_cell[     560] = 32'h9b8adeee;
    ram_cell[     561] = 32'ha61b96bb;
    ram_cell[     562] = 32'hadad985f;
    ram_cell[     563] = 32'haecc01bd;
    ram_cell[     564] = 32'h1ce7849b;
    ram_cell[     565] = 32'h0e276195;
    ram_cell[     566] = 32'h029c9bf7;
    ram_cell[     567] = 32'hb3272d3d;
    ram_cell[     568] = 32'hc9902a9b;
    ram_cell[     569] = 32'h2578d817;
    ram_cell[     570] = 32'h435a8078;
    ram_cell[     571] = 32'h7a387acf;
    ram_cell[     572] = 32'hd8cd6f89;
    ram_cell[     573] = 32'hf5d22c9d;
    ram_cell[     574] = 32'h10b3e878;
    ram_cell[     575] = 32'h1c55dd77;
    ram_cell[     576] = 32'ha9705bff;
    ram_cell[     577] = 32'hdc7a1636;
    ram_cell[     578] = 32'h4535356d;
    ram_cell[     579] = 32'hab1cd975;
    ram_cell[     580] = 32'hcb65f2ba;
    ram_cell[     581] = 32'he52be51a;
    ram_cell[     582] = 32'hf3f0300b;
    ram_cell[     583] = 32'hb33bd9f6;
    ram_cell[     584] = 32'h7d79114b;
    ram_cell[     585] = 32'hf0cedd37;
    ram_cell[     586] = 32'h0450cf1c;
    ram_cell[     587] = 32'hc26fe2fd;
    ram_cell[     588] = 32'hf937ee18;
    ram_cell[     589] = 32'h45bc3da7;
    ram_cell[     590] = 32'hfd667548;
    ram_cell[     591] = 32'h193033b7;
    ram_cell[     592] = 32'he4127aa4;
    ram_cell[     593] = 32'h830a7407;
    ram_cell[     594] = 32'h225fbb15;
    ram_cell[     595] = 32'hfcb9d739;
    ram_cell[     596] = 32'h5b22547b;
    ram_cell[     597] = 32'hc99b259a;
    ram_cell[     598] = 32'hb4a516ee;
    ram_cell[     599] = 32'hcf79fb04;
    ram_cell[     600] = 32'h4d17a0e9;
    ram_cell[     601] = 32'h387b1d6f;
    ram_cell[     602] = 32'hfb9c6378;
    ram_cell[     603] = 32'h0b8b33b6;
    ram_cell[     604] = 32'h3066fd7a;
    ram_cell[     605] = 32'h7047a439;
    ram_cell[     606] = 32'h2cfa72c5;
    ram_cell[     607] = 32'h9582ff02;
    ram_cell[     608] = 32'h3bbc2522;
    ram_cell[     609] = 32'h70c7e1a2;
    ram_cell[     610] = 32'hde56dffb;
    ram_cell[     611] = 32'he81dc09a;
    ram_cell[     612] = 32'h577c7585;
    ram_cell[     613] = 32'hebf3916e;
    ram_cell[     614] = 32'hcd53b909;
    ram_cell[     615] = 32'hf38aa088;
    ram_cell[     616] = 32'h8c93f6b8;
    ram_cell[     617] = 32'h9a65d258;
    ram_cell[     618] = 32'hf3430d38;
    ram_cell[     619] = 32'h7767a0d8;
    ram_cell[     620] = 32'hba4628a8;
    ram_cell[     621] = 32'h13c0141d;
    ram_cell[     622] = 32'h4767ceee;
    ram_cell[     623] = 32'hda06df23;
    ram_cell[     624] = 32'h29598da3;
    ram_cell[     625] = 32'hc3940ceb;
    ram_cell[     626] = 32'ha42e2dc1;
    ram_cell[     627] = 32'h0474a3e5;
    ram_cell[     628] = 32'hb119b68e;
    ram_cell[     629] = 32'h06f3fb9a;
    ram_cell[     630] = 32'hd6df0018;
    ram_cell[     631] = 32'ha2f38818;
    ram_cell[     632] = 32'hacf28c27;
    ram_cell[     633] = 32'ha7394616;
    ram_cell[     634] = 32'h55c70484;
    ram_cell[     635] = 32'hef819b12;
    ram_cell[     636] = 32'h9895db60;
    ram_cell[     637] = 32'h10f13fb1;
    ram_cell[     638] = 32'h6c88530d;
    ram_cell[     639] = 32'h877275ec;
    ram_cell[     640] = 32'h83422a6c;
    ram_cell[     641] = 32'h0b75af1a;
    ram_cell[     642] = 32'hade056a4;
    ram_cell[     643] = 32'hb41ce5ff;
    ram_cell[     644] = 32'h59ee3680;
    ram_cell[     645] = 32'h34e0c478;
    ram_cell[     646] = 32'hbc6f1821;
    ram_cell[     647] = 32'h0dc92375;
    ram_cell[     648] = 32'h2aa95b20;
    ram_cell[     649] = 32'h6f01226f;
    ram_cell[     650] = 32'h32974560;
    ram_cell[     651] = 32'had57c21a;
    ram_cell[     652] = 32'h5feb5ab9;
    ram_cell[     653] = 32'hce504163;
    ram_cell[     654] = 32'h2e3b0510;
    ram_cell[     655] = 32'h6a8199ab;
    ram_cell[     656] = 32'h74f43a92;
    ram_cell[     657] = 32'hed3c13fd;
    ram_cell[     658] = 32'h868dbcc1;
    ram_cell[     659] = 32'h11d3a22c;
    ram_cell[     660] = 32'hf0dc60f6;
    ram_cell[     661] = 32'h2263f8d9;
    ram_cell[     662] = 32'ha604b7c7;
    ram_cell[     663] = 32'h32d0a7f4;
    ram_cell[     664] = 32'h33c0226f;
    ram_cell[     665] = 32'hff0402fa;
    ram_cell[     666] = 32'h51d7a4c6;
    ram_cell[     667] = 32'h0755f9b7;
    ram_cell[     668] = 32'h7d474157;
    ram_cell[     669] = 32'heedc7f7d;
    ram_cell[     670] = 32'hf799b09a;
    ram_cell[     671] = 32'h798cbe15;
    ram_cell[     672] = 32'hc3e6c4f0;
    ram_cell[     673] = 32'h5cb089e3;
    ram_cell[     674] = 32'hd1546c15;
    ram_cell[     675] = 32'h30999e68;
    ram_cell[     676] = 32'h1fe26353;
    ram_cell[     677] = 32'h890bee5e;
    ram_cell[     678] = 32'h74a0810d;
    ram_cell[     679] = 32'h5e906ab1;
    ram_cell[     680] = 32'ha800d3c4;
    ram_cell[     681] = 32'h295e7cf6;
    ram_cell[     682] = 32'hac64b09b;
    ram_cell[     683] = 32'hf935b581;
    ram_cell[     684] = 32'h700c0bb0;
    ram_cell[     685] = 32'hf24b219b;
    ram_cell[     686] = 32'h14306340;
    ram_cell[     687] = 32'h8d0b1a49;
    ram_cell[     688] = 32'h7bc49d53;
    ram_cell[     689] = 32'h9d851bc5;
    ram_cell[     690] = 32'he9cbf748;
    ram_cell[     691] = 32'hf1c77034;
    ram_cell[     692] = 32'hd5e97faf;
    ram_cell[     693] = 32'h0ceaad4e;
    ram_cell[     694] = 32'h31c455ac;
    ram_cell[     695] = 32'h12ec6909;
    ram_cell[     696] = 32'h35a78220;
    ram_cell[     697] = 32'h32647519;
    ram_cell[     698] = 32'h2a0e2fa0;
    ram_cell[     699] = 32'hfaaf107b;
    ram_cell[     700] = 32'hba3b4036;
    ram_cell[     701] = 32'hd533830f;
    ram_cell[     702] = 32'h61c54dc3;
    ram_cell[     703] = 32'h59b62089;
    ram_cell[     704] = 32'h9c60aae2;
    ram_cell[     705] = 32'h41142ffa;
    ram_cell[     706] = 32'h9dd6905c;
    ram_cell[     707] = 32'he0564bd9;
    ram_cell[     708] = 32'hf6cf9c4f;
    ram_cell[     709] = 32'hdfad2504;
    ram_cell[     710] = 32'h7c1d62a2;
    ram_cell[     711] = 32'h92bac1eb;
    ram_cell[     712] = 32'ha40babf5;
    ram_cell[     713] = 32'hbfcbc3ea;
    ram_cell[     714] = 32'hbbc0ab3e;
    ram_cell[     715] = 32'h31877d51;
    ram_cell[     716] = 32'hcd983518;
    ram_cell[     717] = 32'h8f5d3b30;
    ram_cell[     718] = 32'h8b6ca075;
    ram_cell[     719] = 32'h69a4efc8;
    ram_cell[     720] = 32'he7bde55c;
    ram_cell[     721] = 32'h64e8248d;
    ram_cell[     722] = 32'h78f39722;
    ram_cell[     723] = 32'h58612128;
    ram_cell[     724] = 32'h3b99eb58;
    ram_cell[     725] = 32'hd40e8b5b;
    ram_cell[     726] = 32'h93129202;
    ram_cell[     727] = 32'h6f6303ab;
    ram_cell[     728] = 32'hf8471349;
    ram_cell[     729] = 32'h39fc86ea;
    ram_cell[     730] = 32'h8fa7486f;
    ram_cell[     731] = 32'hcab1186f;
    ram_cell[     732] = 32'h654e4394;
    ram_cell[     733] = 32'h6fdf4138;
    ram_cell[     734] = 32'h6730768c;
    ram_cell[     735] = 32'hae80e12d;
    ram_cell[     736] = 32'hcaf9d45a;
    ram_cell[     737] = 32'hfddb04b2;
    ram_cell[     738] = 32'h3a493326;
    ram_cell[     739] = 32'h04866315;
    ram_cell[     740] = 32'h8de0b6fa;
    ram_cell[     741] = 32'h539ac9d1;
    ram_cell[     742] = 32'h2819fd4a;
    ram_cell[     743] = 32'h5f9c3d8b;
    ram_cell[     744] = 32'hc9693c10;
    ram_cell[     745] = 32'hdccdf8c7;
    ram_cell[     746] = 32'h0344d29f;
    ram_cell[     747] = 32'h16659d11;
    ram_cell[     748] = 32'hd84a61c9;
    ram_cell[     749] = 32'h07318046;
    ram_cell[     750] = 32'hb01a1aca;
    ram_cell[     751] = 32'h633bcc31;
    ram_cell[     752] = 32'hd291e56e;
    ram_cell[     753] = 32'h69e15fee;
    ram_cell[     754] = 32'h236287e7;
    ram_cell[     755] = 32'h195afafc;
    ram_cell[     756] = 32'hdfa42f81;
    ram_cell[     757] = 32'h8146cc86;
    ram_cell[     758] = 32'h4f9054bc;
    ram_cell[     759] = 32'hd078a4e4;
    ram_cell[     760] = 32'h98ae4165;
    ram_cell[     761] = 32'hbb71cd47;
    ram_cell[     762] = 32'h7596984c;
    ram_cell[     763] = 32'hb197bd86;
    ram_cell[     764] = 32'hdc315356;
    ram_cell[     765] = 32'he0c181db;
    ram_cell[     766] = 32'h8959d67d;
    ram_cell[     767] = 32'h381d509f;
end

endmodule

