
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hdbb421a4;
    ram_cell[       1] = 32'h0;  // 32'hcac16870;
    ram_cell[       2] = 32'h0;  // 32'h5ebd1d54;
    ram_cell[       3] = 32'h0;  // 32'h25ce31e1;
    ram_cell[       4] = 32'h0;  // 32'hdb01f2a0;
    ram_cell[       5] = 32'h0;  // 32'he9477bfe;
    ram_cell[       6] = 32'h0;  // 32'h2473210f;
    ram_cell[       7] = 32'h0;  // 32'h0da0e4e8;
    ram_cell[       8] = 32'h0;  // 32'h4c1f3af7;
    ram_cell[       9] = 32'h0;  // 32'hdf6da0b2;
    ram_cell[      10] = 32'h0;  // 32'hc4d24154;
    ram_cell[      11] = 32'h0;  // 32'h624d390a;
    ram_cell[      12] = 32'h0;  // 32'h3a1097e0;
    ram_cell[      13] = 32'h0;  // 32'h779b01b6;
    ram_cell[      14] = 32'h0;  // 32'h01a0ce64;
    ram_cell[      15] = 32'h0;  // 32'hf3e0e017;
    ram_cell[      16] = 32'h0;  // 32'heabbdf55;
    ram_cell[      17] = 32'h0;  // 32'hfd1b2971;
    ram_cell[      18] = 32'h0;  // 32'h67d0eaef;
    ram_cell[      19] = 32'h0;  // 32'hb47c5e57;
    ram_cell[      20] = 32'h0;  // 32'h7923d19d;
    ram_cell[      21] = 32'h0;  // 32'h64fbb3b9;
    ram_cell[      22] = 32'h0;  // 32'h93019c7d;
    ram_cell[      23] = 32'h0;  // 32'h10e3b519;
    ram_cell[      24] = 32'h0;  // 32'hed25b2a0;
    ram_cell[      25] = 32'h0;  // 32'hbd5c197f;
    ram_cell[      26] = 32'h0;  // 32'hec253af2;
    ram_cell[      27] = 32'h0;  // 32'hcb061767;
    ram_cell[      28] = 32'h0;  // 32'hac7834bc;
    ram_cell[      29] = 32'h0;  // 32'h7e004ca7;
    ram_cell[      30] = 32'h0;  // 32'hc0c56539;
    ram_cell[      31] = 32'h0;  // 32'h90b394c5;
    ram_cell[      32] = 32'h0;  // 32'h6b8235c9;
    ram_cell[      33] = 32'h0;  // 32'h05e855aa;
    ram_cell[      34] = 32'h0;  // 32'hd41961af;
    ram_cell[      35] = 32'h0;  // 32'hbae3c16d;
    ram_cell[      36] = 32'h0;  // 32'hae0bc92b;
    ram_cell[      37] = 32'h0;  // 32'h29ef4b00;
    ram_cell[      38] = 32'h0;  // 32'heee4e742;
    ram_cell[      39] = 32'h0;  // 32'h19f3e9e1;
    ram_cell[      40] = 32'h0;  // 32'h00230f9a;
    ram_cell[      41] = 32'h0;  // 32'h77c335dc;
    ram_cell[      42] = 32'h0;  // 32'hce427823;
    ram_cell[      43] = 32'h0;  // 32'h6bff84ce;
    ram_cell[      44] = 32'h0;  // 32'hc1b5653a;
    ram_cell[      45] = 32'h0;  // 32'hbbcf5be7;
    ram_cell[      46] = 32'h0;  // 32'hcd98766a;
    ram_cell[      47] = 32'h0;  // 32'he07efdfe;
    ram_cell[      48] = 32'h0;  // 32'h39a2383e;
    ram_cell[      49] = 32'h0;  // 32'hee1c7a7d;
    ram_cell[      50] = 32'h0;  // 32'hd1ccbd50;
    ram_cell[      51] = 32'h0;  // 32'h6b7f445e;
    ram_cell[      52] = 32'h0;  // 32'hdb207acd;
    ram_cell[      53] = 32'h0;  // 32'hcae40621;
    ram_cell[      54] = 32'h0;  // 32'he9b5a4dd;
    ram_cell[      55] = 32'h0;  // 32'h49929cb5;
    ram_cell[      56] = 32'h0;  // 32'h45ab897c;
    ram_cell[      57] = 32'h0;  // 32'h14167907;
    ram_cell[      58] = 32'h0;  // 32'h7bb87d76;
    ram_cell[      59] = 32'h0;  // 32'hc4571163;
    ram_cell[      60] = 32'h0;  // 32'h27d9345c;
    ram_cell[      61] = 32'h0;  // 32'h15008b78;
    ram_cell[      62] = 32'h0;  // 32'hfa46d0fc;
    ram_cell[      63] = 32'h0;  // 32'hffb1b6be;
    ram_cell[      64] = 32'h0;  // 32'hbd4bd689;
    ram_cell[      65] = 32'h0;  // 32'hbfce9aff;
    ram_cell[      66] = 32'h0;  // 32'hceedc18a;
    ram_cell[      67] = 32'h0;  // 32'h359e6c15;
    ram_cell[      68] = 32'h0;  // 32'h0d0e7aaf;
    ram_cell[      69] = 32'h0;  // 32'h333894d8;
    ram_cell[      70] = 32'h0;  // 32'he8b5e180;
    ram_cell[      71] = 32'h0;  // 32'h311f21e4;
    ram_cell[      72] = 32'h0;  // 32'h73713b66;
    ram_cell[      73] = 32'h0;  // 32'h161274bf;
    ram_cell[      74] = 32'h0;  // 32'hbd193867;
    ram_cell[      75] = 32'h0;  // 32'h7a7dfcf6;
    ram_cell[      76] = 32'h0;  // 32'hc6f283ad;
    ram_cell[      77] = 32'h0;  // 32'h7b2a3170;
    ram_cell[      78] = 32'h0;  // 32'h946ce8e0;
    ram_cell[      79] = 32'h0;  // 32'hca63fa60;
    ram_cell[      80] = 32'h0;  // 32'ha092ef57;
    ram_cell[      81] = 32'h0;  // 32'hc6dddd9a;
    ram_cell[      82] = 32'h0;  // 32'h971fd29f;
    ram_cell[      83] = 32'h0;  // 32'h4cd4a0ac;
    ram_cell[      84] = 32'h0;  // 32'h0dcdd589;
    ram_cell[      85] = 32'h0;  // 32'h8fac8679;
    ram_cell[      86] = 32'h0;  // 32'ha23001e1;
    ram_cell[      87] = 32'h0;  // 32'hc4debdcf;
    ram_cell[      88] = 32'h0;  // 32'h5832d33d;
    ram_cell[      89] = 32'h0;  // 32'h1831e9e0;
    ram_cell[      90] = 32'h0;  // 32'h7d18a40b;
    ram_cell[      91] = 32'h0;  // 32'hdf2135b2;
    ram_cell[      92] = 32'h0;  // 32'h40a1b169;
    ram_cell[      93] = 32'h0;  // 32'haf7958cc;
    ram_cell[      94] = 32'h0;  // 32'h6ea66c01;
    ram_cell[      95] = 32'h0;  // 32'hb5c3e353;
    ram_cell[      96] = 32'h0;  // 32'h8c19bb8f;
    ram_cell[      97] = 32'h0;  // 32'h26281f6f;
    ram_cell[      98] = 32'h0;  // 32'hc234939f;
    ram_cell[      99] = 32'h0;  // 32'h1a7c3699;
    ram_cell[     100] = 32'h0;  // 32'hbf9927cd;
    ram_cell[     101] = 32'h0;  // 32'hd097f9e8;
    ram_cell[     102] = 32'h0;  // 32'h74002e14;
    ram_cell[     103] = 32'h0;  // 32'he7f6d672;
    ram_cell[     104] = 32'h0;  // 32'h073e92bf;
    ram_cell[     105] = 32'h0;  // 32'hdfed6a77;
    ram_cell[     106] = 32'h0;  // 32'h66abb665;
    ram_cell[     107] = 32'h0;  // 32'h0897e958;
    ram_cell[     108] = 32'h0;  // 32'h826efc2e;
    ram_cell[     109] = 32'h0;  // 32'hc3676ed5;
    ram_cell[     110] = 32'h0;  // 32'hbca0aa54;
    ram_cell[     111] = 32'h0;  // 32'h51cc7d58;
    ram_cell[     112] = 32'h0;  // 32'hd00f1bc3;
    ram_cell[     113] = 32'h0;  // 32'h6bd05990;
    ram_cell[     114] = 32'h0;  // 32'hde3d271a;
    ram_cell[     115] = 32'h0;  // 32'hb98747a8;
    ram_cell[     116] = 32'h0;  // 32'h48cc1159;
    ram_cell[     117] = 32'h0;  // 32'hc58a6bb5;
    ram_cell[     118] = 32'h0;  // 32'hc3b752dc;
    ram_cell[     119] = 32'h0;  // 32'hf8cd1d6a;
    ram_cell[     120] = 32'h0;  // 32'h836b803d;
    ram_cell[     121] = 32'h0;  // 32'h89f4c930;
    ram_cell[     122] = 32'h0;  // 32'h5d32970a;
    ram_cell[     123] = 32'h0;  // 32'h9bf56a67;
    ram_cell[     124] = 32'h0;  // 32'hd4d56256;
    ram_cell[     125] = 32'h0;  // 32'h7d60ddcb;
    ram_cell[     126] = 32'h0;  // 32'h9b360470;
    ram_cell[     127] = 32'h0;  // 32'hf571fa87;
    ram_cell[     128] = 32'h0;  // 32'h7bc8d6ca;
    ram_cell[     129] = 32'h0;  // 32'hf2b9d17b;
    ram_cell[     130] = 32'h0;  // 32'h717e2ff0;
    ram_cell[     131] = 32'h0;  // 32'ha14d1f57;
    ram_cell[     132] = 32'h0;  // 32'h5c9b3646;
    ram_cell[     133] = 32'h0;  // 32'h04b8c244;
    ram_cell[     134] = 32'h0;  // 32'h8a14792f;
    ram_cell[     135] = 32'h0;  // 32'h9882229f;
    ram_cell[     136] = 32'h0;  // 32'hb81e2889;
    ram_cell[     137] = 32'h0;  // 32'h7f73e7c4;
    ram_cell[     138] = 32'h0;  // 32'h0e679a93;
    ram_cell[     139] = 32'h0;  // 32'h17c62f37;
    ram_cell[     140] = 32'h0;  // 32'hb74cc18e;
    ram_cell[     141] = 32'h0;  // 32'haf6006e7;
    ram_cell[     142] = 32'h0;  // 32'h0b895fa5;
    ram_cell[     143] = 32'h0;  // 32'h9b39c91e;
    ram_cell[     144] = 32'h0;  // 32'h83ce8885;
    ram_cell[     145] = 32'h0;  // 32'hc105a489;
    ram_cell[     146] = 32'h0;  // 32'h79bd2484;
    ram_cell[     147] = 32'h0;  // 32'hd3f86b40;
    ram_cell[     148] = 32'h0;  // 32'ha318684f;
    ram_cell[     149] = 32'h0;  // 32'hdaf3fafc;
    ram_cell[     150] = 32'h0;  // 32'h2128a2d9;
    ram_cell[     151] = 32'h0;  // 32'h2f6f3c64;
    ram_cell[     152] = 32'h0;  // 32'hb8742d75;
    ram_cell[     153] = 32'h0;  // 32'hcc2bd3d5;
    ram_cell[     154] = 32'h0;  // 32'h547dda4e;
    ram_cell[     155] = 32'h0;  // 32'hf4620163;
    ram_cell[     156] = 32'h0;  // 32'h22a82a81;
    ram_cell[     157] = 32'h0;  // 32'he7d7a844;
    ram_cell[     158] = 32'h0;  // 32'h02db6749;
    ram_cell[     159] = 32'h0;  // 32'h6ca7ef33;
    ram_cell[     160] = 32'h0;  // 32'he2bc3834;
    ram_cell[     161] = 32'h0;  // 32'h607eff56;
    ram_cell[     162] = 32'h0;  // 32'h708427ee;
    ram_cell[     163] = 32'h0;  // 32'h0235899e;
    ram_cell[     164] = 32'h0;  // 32'h1fef689c;
    ram_cell[     165] = 32'h0;  // 32'h59029420;
    ram_cell[     166] = 32'h0;  // 32'hc524bb9a;
    ram_cell[     167] = 32'h0;  // 32'hbf53b9af;
    ram_cell[     168] = 32'h0;  // 32'h1be9ca5c;
    ram_cell[     169] = 32'h0;  // 32'h78832458;
    ram_cell[     170] = 32'h0;  // 32'h0a591a2e;
    ram_cell[     171] = 32'h0;  // 32'h8e31fe12;
    ram_cell[     172] = 32'h0;  // 32'h337981e5;
    ram_cell[     173] = 32'h0;  // 32'haa5af660;
    ram_cell[     174] = 32'h0;  // 32'h15936611;
    ram_cell[     175] = 32'h0;  // 32'h87acef75;
    ram_cell[     176] = 32'h0;  // 32'h539e1785;
    ram_cell[     177] = 32'h0;  // 32'h9e3197a6;
    ram_cell[     178] = 32'h0;  // 32'h276a93ac;
    ram_cell[     179] = 32'h0;  // 32'h92b68fe9;
    ram_cell[     180] = 32'h0;  // 32'h8d7e6aaa;
    ram_cell[     181] = 32'h0;  // 32'hb40c039a;
    ram_cell[     182] = 32'h0;  // 32'hc426a255;
    ram_cell[     183] = 32'h0;  // 32'h01efddb5;
    ram_cell[     184] = 32'h0;  // 32'h66f58c8a;
    ram_cell[     185] = 32'h0;  // 32'h140436ce;
    ram_cell[     186] = 32'h0;  // 32'h66dc0353;
    ram_cell[     187] = 32'h0;  // 32'h669e98e8;
    ram_cell[     188] = 32'h0;  // 32'h7c76c2d0;
    ram_cell[     189] = 32'h0;  // 32'ha8c8a7ad;
    ram_cell[     190] = 32'h0;  // 32'h731cefc5;
    ram_cell[     191] = 32'h0;  // 32'ha12cbb83;
    ram_cell[     192] = 32'h0;  // 32'h66366bee;
    ram_cell[     193] = 32'h0;  // 32'h1ffeda9f;
    ram_cell[     194] = 32'h0;  // 32'h3d209ca8;
    ram_cell[     195] = 32'h0;  // 32'hb972855e;
    ram_cell[     196] = 32'h0;  // 32'hb3cb8473;
    ram_cell[     197] = 32'h0;  // 32'h2e4c7e49;
    ram_cell[     198] = 32'h0;  // 32'hb823c36a;
    ram_cell[     199] = 32'h0;  // 32'h2e7d13c1;
    ram_cell[     200] = 32'h0;  // 32'h4bab3467;
    ram_cell[     201] = 32'h0;  // 32'hd65f952e;
    ram_cell[     202] = 32'h0;  // 32'h523d44da;
    ram_cell[     203] = 32'h0;  // 32'h817148f5;
    ram_cell[     204] = 32'h0;  // 32'h010f03c8;
    ram_cell[     205] = 32'h0;  // 32'h1d4db6e5;
    ram_cell[     206] = 32'h0;  // 32'h81478a9d;
    ram_cell[     207] = 32'h0;  // 32'h7badfbe1;
    ram_cell[     208] = 32'h0;  // 32'h2fdeadcb;
    ram_cell[     209] = 32'h0;  // 32'h4cd7d3f3;
    ram_cell[     210] = 32'h0;  // 32'hb65b4b67;
    ram_cell[     211] = 32'h0;  // 32'h54f627c6;
    ram_cell[     212] = 32'h0;  // 32'hf0aedfd8;
    ram_cell[     213] = 32'h0;  // 32'h61cd27f3;
    ram_cell[     214] = 32'h0;  // 32'h4229294b;
    ram_cell[     215] = 32'h0;  // 32'h840580f8;
    ram_cell[     216] = 32'h0;  // 32'h68801817;
    ram_cell[     217] = 32'h0;  // 32'hbc3f24d5;
    ram_cell[     218] = 32'h0;  // 32'h28611f9a;
    ram_cell[     219] = 32'h0;  // 32'h5f96e81a;
    ram_cell[     220] = 32'h0;  // 32'hbffb2c4a;
    ram_cell[     221] = 32'h0;  // 32'hc69a0b85;
    ram_cell[     222] = 32'h0;  // 32'h93968019;
    ram_cell[     223] = 32'h0;  // 32'h89972754;
    ram_cell[     224] = 32'h0;  // 32'he4e6382d;
    ram_cell[     225] = 32'h0;  // 32'hb3fae818;
    ram_cell[     226] = 32'h0;  // 32'h4af8c179;
    ram_cell[     227] = 32'h0;  // 32'hdf7e2bab;
    ram_cell[     228] = 32'h0;  // 32'h57eccdc8;
    ram_cell[     229] = 32'h0;  // 32'h0977ba3d;
    ram_cell[     230] = 32'h0;  // 32'hf7743342;
    ram_cell[     231] = 32'h0;  // 32'h94896f9a;
    ram_cell[     232] = 32'h0;  // 32'h596a0d98;
    ram_cell[     233] = 32'h0;  // 32'h23efef73;
    ram_cell[     234] = 32'h0;  // 32'h3bdd76cd;
    ram_cell[     235] = 32'h0;  // 32'h9fa0c6ee;
    ram_cell[     236] = 32'h0;  // 32'h6d03f550;
    ram_cell[     237] = 32'h0;  // 32'hfc00fdc9;
    ram_cell[     238] = 32'h0;  // 32'h13c349c5;
    ram_cell[     239] = 32'h0;  // 32'h6b84afc7;
    ram_cell[     240] = 32'h0;  // 32'h89f935b8;
    ram_cell[     241] = 32'h0;  // 32'hd216b4c4;
    ram_cell[     242] = 32'h0;  // 32'hae8198a9;
    ram_cell[     243] = 32'h0;  // 32'hb0e3c9d5;
    ram_cell[     244] = 32'h0;  // 32'h89f86004;
    ram_cell[     245] = 32'h0;  // 32'h6f62dcc5;
    ram_cell[     246] = 32'h0;  // 32'hf6647d78;
    ram_cell[     247] = 32'h0;  // 32'h521a1bb1;
    ram_cell[     248] = 32'h0;  // 32'h3b22c81d;
    ram_cell[     249] = 32'h0;  // 32'haf8661d3;
    ram_cell[     250] = 32'h0;  // 32'hecf0d8e2;
    ram_cell[     251] = 32'h0;  // 32'hc281117e;
    ram_cell[     252] = 32'h0;  // 32'h745d1f15;
    ram_cell[     253] = 32'h0;  // 32'hcdc67203;
    ram_cell[     254] = 32'h0;  // 32'h94775c20;
    ram_cell[     255] = 32'h0;  // 32'h81a2ad86;
    // src matrix A
    ram_cell[     256] = 32'hf784f3be;
    ram_cell[     257] = 32'hde258d52;
    ram_cell[     258] = 32'h6bdee95a;
    ram_cell[     259] = 32'h29b8f94b;
    ram_cell[     260] = 32'h7838aa93;
    ram_cell[     261] = 32'hedfef778;
    ram_cell[     262] = 32'h59f91f7d;
    ram_cell[     263] = 32'h2921a8a2;
    ram_cell[     264] = 32'h05427b72;
    ram_cell[     265] = 32'h673cdfe5;
    ram_cell[     266] = 32'h97b983fc;
    ram_cell[     267] = 32'h36416fa4;
    ram_cell[     268] = 32'he71c8a41;
    ram_cell[     269] = 32'h3526f230;
    ram_cell[     270] = 32'h3a0558ec;
    ram_cell[     271] = 32'h47630449;
    ram_cell[     272] = 32'h3aba979d;
    ram_cell[     273] = 32'hfa7aa0d9;
    ram_cell[     274] = 32'hba02861e;
    ram_cell[     275] = 32'h49457773;
    ram_cell[     276] = 32'h88f96e8a;
    ram_cell[     277] = 32'h01a307a4;
    ram_cell[     278] = 32'h7eab406e;
    ram_cell[     279] = 32'h2dd0666f;
    ram_cell[     280] = 32'hadb6ecbf;
    ram_cell[     281] = 32'h586c2e72;
    ram_cell[     282] = 32'hdfbf3af3;
    ram_cell[     283] = 32'h32ef3b29;
    ram_cell[     284] = 32'h88b1fb6c;
    ram_cell[     285] = 32'h58f5d0d4;
    ram_cell[     286] = 32'hf59c8c6d;
    ram_cell[     287] = 32'h335078b5;
    ram_cell[     288] = 32'h78f532c1;
    ram_cell[     289] = 32'h0ca4728d;
    ram_cell[     290] = 32'hc6cd6c15;
    ram_cell[     291] = 32'hd9d1c7a4;
    ram_cell[     292] = 32'h4c60c586;
    ram_cell[     293] = 32'h95dd4214;
    ram_cell[     294] = 32'h050fa313;
    ram_cell[     295] = 32'hb9ebbd8b;
    ram_cell[     296] = 32'hab079a04;
    ram_cell[     297] = 32'hf25920f4;
    ram_cell[     298] = 32'hb20f1f2d;
    ram_cell[     299] = 32'h30226ae1;
    ram_cell[     300] = 32'hc89dc5d2;
    ram_cell[     301] = 32'h2513966b;
    ram_cell[     302] = 32'h74ca5131;
    ram_cell[     303] = 32'h303cba1c;
    ram_cell[     304] = 32'h8d2f7d0b;
    ram_cell[     305] = 32'h80d2397a;
    ram_cell[     306] = 32'heb892b5f;
    ram_cell[     307] = 32'ha72b3fa6;
    ram_cell[     308] = 32'h86bc2bf5;
    ram_cell[     309] = 32'hdbdbcd29;
    ram_cell[     310] = 32'h46b62f17;
    ram_cell[     311] = 32'h70f11287;
    ram_cell[     312] = 32'hd6a3ac48;
    ram_cell[     313] = 32'h8bc807cc;
    ram_cell[     314] = 32'h19c8e62f;
    ram_cell[     315] = 32'h93c24f3e;
    ram_cell[     316] = 32'h0dfde43c;
    ram_cell[     317] = 32'h562ae742;
    ram_cell[     318] = 32'h1265aed8;
    ram_cell[     319] = 32'h9809e570;
    ram_cell[     320] = 32'hd836ce77;
    ram_cell[     321] = 32'hbfb865b4;
    ram_cell[     322] = 32'h8169fda6;
    ram_cell[     323] = 32'h519ee9cc;
    ram_cell[     324] = 32'hd755d1fe;
    ram_cell[     325] = 32'h3c0e4a86;
    ram_cell[     326] = 32'hff984c82;
    ram_cell[     327] = 32'hc6af3142;
    ram_cell[     328] = 32'h8b85b0f3;
    ram_cell[     329] = 32'h432666d0;
    ram_cell[     330] = 32'h342d1bc0;
    ram_cell[     331] = 32'h11cc2265;
    ram_cell[     332] = 32'h37d738ee;
    ram_cell[     333] = 32'hfc598f94;
    ram_cell[     334] = 32'hdde1cf51;
    ram_cell[     335] = 32'hb5eda7a9;
    ram_cell[     336] = 32'hc3a45f77;
    ram_cell[     337] = 32'h78e57549;
    ram_cell[     338] = 32'heaeb9e01;
    ram_cell[     339] = 32'h546bf634;
    ram_cell[     340] = 32'hf202cda1;
    ram_cell[     341] = 32'h7fe4c165;
    ram_cell[     342] = 32'h0dddd585;
    ram_cell[     343] = 32'h05f3893b;
    ram_cell[     344] = 32'ha8de0c2a;
    ram_cell[     345] = 32'h321412d5;
    ram_cell[     346] = 32'h2cb61c6d;
    ram_cell[     347] = 32'h849bb858;
    ram_cell[     348] = 32'h77a8561e;
    ram_cell[     349] = 32'h8893ab69;
    ram_cell[     350] = 32'hb5cdb53e;
    ram_cell[     351] = 32'h904ce0fa;
    ram_cell[     352] = 32'h20a5dfd1;
    ram_cell[     353] = 32'h44bda8e6;
    ram_cell[     354] = 32'h33c61bcc;
    ram_cell[     355] = 32'ha58404e6;
    ram_cell[     356] = 32'h1a86528c;
    ram_cell[     357] = 32'h9d8cd9d1;
    ram_cell[     358] = 32'hfde3db18;
    ram_cell[     359] = 32'hd2ae4204;
    ram_cell[     360] = 32'h0a3fc2cc;
    ram_cell[     361] = 32'h567f3c54;
    ram_cell[     362] = 32'h5882f549;
    ram_cell[     363] = 32'h2476bec1;
    ram_cell[     364] = 32'h33b71b8c;
    ram_cell[     365] = 32'hf96343af;
    ram_cell[     366] = 32'h86f6f1b8;
    ram_cell[     367] = 32'h53c0103e;
    ram_cell[     368] = 32'hac8081d3;
    ram_cell[     369] = 32'h98e61c86;
    ram_cell[     370] = 32'hf1292a77;
    ram_cell[     371] = 32'h8e42d2e8;
    ram_cell[     372] = 32'h0b98a871;
    ram_cell[     373] = 32'h281f4a74;
    ram_cell[     374] = 32'h0cb535ba;
    ram_cell[     375] = 32'hfac1f448;
    ram_cell[     376] = 32'hd73113c9;
    ram_cell[     377] = 32'h152a59e6;
    ram_cell[     378] = 32'h55ca6bbd;
    ram_cell[     379] = 32'hf2483e4c;
    ram_cell[     380] = 32'hde5c59e6;
    ram_cell[     381] = 32'h83e22eb5;
    ram_cell[     382] = 32'h4b848eee;
    ram_cell[     383] = 32'ha3abbec7;
    ram_cell[     384] = 32'h48b6ebf7;
    ram_cell[     385] = 32'h09cf523f;
    ram_cell[     386] = 32'h18f227d2;
    ram_cell[     387] = 32'h0cf62d85;
    ram_cell[     388] = 32'hac9f6e88;
    ram_cell[     389] = 32'hcb1a35a6;
    ram_cell[     390] = 32'hf6f6c6a7;
    ram_cell[     391] = 32'h9e2c2644;
    ram_cell[     392] = 32'h66828a2c;
    ram_cell[     393] = 32'hb84b02a3;
    ram_cell[     394] = 32'hd61a1661;
    ram_cell[     395] = 32'h12c0702b;
    ram_cell[     396] = 32'h0cda7548;
    ram_cell[     397] = 32'h4b1eb18e;
    ram_cell[     398] = 32'h2949dfd0;
    ram_cell[     399] = 32'h985e2119;
    ram_cell[     400] = 32'h22873a6b;
    ram_cell[     401] = 32'h0b2221f0;
    ram_cell[     402] = 32'he2ee38ae;
    ram_cell[     403] = 32'h4c2a3fa5;
    ram_cell[     404] = 32'h5241775e;
    ram_cell[     405] = 32'h092acbb4;
    ram_cell[     406] = 32'h951cf1b8;
    ram_cell[     407] = 32'h0d59062c;
    ram_cell[     408] = 32'h15af4cc8;
    ram_cell[     409] = 32'h09831d41;
    ram_cell[     410] = 32'h1d6527db;
    ram_cell[     411] = 32'h7d2cb29e;
    ram_cell[     412] = 32'h1ae566f1;
    ram_cell[     413] = 32'hd87dce33;
    ram_cell[     414] = 32'hed0e44a3;
    ram_cell[     415] = 32'h59565a0e;
    ram_cell[     416] = 32'h7db903da;
    ram_cell[     417] = 32'h2a0c2881;
    ram_cell[     418] = 32'h553fc54f;
    ram_cell[     419] = 32'h1ddc4edb;
    ram_cell[     420] = 32'h9fa7719a;
    ram_cell[     421] = 32'h9a073691;
    ram_cell[     422] = 32'h53e2bc2a;
    ram_cell[     423] = 32'h8a67ca84;
    ram_cell[     424] = 32'hac84521f;
    ram_cell[     425] = 32'h7ea120ed;
    ram_cell[     426] = 32'h5844225c;
    ram_cell[     427] = 32'hc18ade7f;
    ram_cell[     428] = 32'hc48efa53;
    ram_cell[     429] = 32'h46248f7a;
    ram_cell[     430] = 32'heed902a0;
    ram_cell[     431] = 32'h48886807;
    ram_cell[     432] = 32'h848abd95;
    ram_cell[     433] = 32'h6997745f;
    ram_cell[     434] = 32'h06e48106;
    ram_cell[     435] = 32'h210e25e0;
    ram_cell[     436] = 32'h4a440b58;
    ram_cell[     437] = 32'hc1f06067;
    ram_cell[     438] = 32'h23b1737c;
    ram_cell[     439] = 32'h50a7a2b4;
    ram_cell[     440] = 32'h7f51c809;
    ram_cell[     441] = 32'h9827f826;
    ram_cell[     442] = 32'h84835472;
    ram_cell[     443] = 32'h2b7f2d2d;
    ram_cell[     444] = 32'h484ca937;
    ram_cell[     445] = 32'h97719f4b;
    ram_cell[     446] = 32'h82d21925;
    ram_cell[     447] = 32'h7a468ae2;
    ram_cell[     448] = 32'hd2d06bb7;
    ram_cell[     449] = 32'h507053f7;
    ram_cell[     450] = 32'h114e07da;
    ram_cell[     451] = 32'h95f18117;
    ram_cell[     452] = 32'h1fc56f76;
    ram_cell[     453] = 32'he8e785fa;
    ram_cell[     454] = 32'hb8802ee2;
    ram_cell[     455] = 32'hbfbd68d9;
    ram_cell[     456] = 32'h54fa6757;
    ram_cell[     457] = 32'h6fd573d0;
    ram_cell[     458] = 32'h0f93aa6f;
    ram_cell[     459] = 32'ha04561c7;
    ram_cell[     460] = 32'h1deb29b0;
    ram_cell[     461] = 32'he7a6ebff;
    ram_cell[     462] = 32'h863dcf36;
    ram_cell[     463] = 32'ha0dd101a;
    ram_cell[     464] = 32'h5f43d65b;
    ram_cell[     465] = 32'h743384e1;
    ram_cell[     466] = 32'hcf615271;
    ram_cell[     467] = 32'h8c8abbdb;
    ram_cell[     468] = 32'hed1fe879;
    ram_cell[     469] = 32'h90716b32;
    ram_cell[     470] = 32'h2e86bf65;
    ram_cell[     471] = 32'h660dc473;
    ram_cell[     472] = 32'hfa058023;
    ram_cell[     473] = 32'h15b23878;
    ram_cell[     474] = 32'ha7514c14;
    ram_cell[     475] = 32'h854f1a52;
    ram_cell[     476] = 32'h45fc266a;
    ram_cell[     477] = 32'h105e3262;
    ram_cell[     478] = 32'h5854081a;
    ram_cell[     479] = 32'h630693ee;
    ram_cell[     480] = 32'ha4de56ba;
    ram_cell[     481] = 32'he6d1d268;
    ram_cell[     482] = 32'h0bc4bdb1;
    ram_cell[     483] = 32'h617c037d;
    ram_cell[     484] = 32'h2f788732;
    ram_cell[     485] = 32'he97a3be3;
    ram_cell[     486] = 32'hae1a09a0;
    ram_cell[     487] = 32'h55045dc2;
    ram_cell[     488] = 32'h25094ded;
    ram_cell[     489] = 32'h72abd00d;
    ram_cell[     490] = 32'h99d16494;
    ram_cell[     491] = 32'h13086e73;
    ram_cell[     492] = 32'hd0d72da8;
    ram_cell[     493] = 32'hc86beb3b;
    ram_cell[     494] = 32'hb9a92557;
    ram_cell[     495] = 32'hf79a663e;
    ram_cell[     496] = 32'hd8ea3e60;
    ram_cell[     497] = 32'h1cf6c9c5;
    ram_cell[     498] = 32'heac65dab;
    ram_cell[     499] = 32'he92e06ab;
    ram_cell[     500] = 32'h95262789;
    ram_cell[     501] = 32'h049fa9cf;
    ram_cell[     502] = 32'h226f6e4f;
    ram_cell[     503] = 32'hff75b1c4;
    ram_cell[     504] = 32'hc9cef19b;
    ram_cell[     505] = 32'he6ff9279;
    ram_cell[     506] = 32'h79e7b742;
    ram_cell[     507] = 32'h64d7039c;
    ram_cell[     508] = 32'h60cfcc89;
    ram_cell[     509] = 32'h221f5532;
    ram_cell[     510] = 32'h5e2a9e88;
    ram_cell[     511] = 32'hb5b081e9;
    // src matrix B
    ram_cell[     512] = 32'ha791a39d;
    ram_cell[     513] = 32'h97a5fb42;
    ram_cell[     514] = 32'hd17a977d;
    ram_cell[     515] = 32'h2818283a;
    ram_cell[     516] = 32'h5b067f9e;
    ram_cell[     517] = 32'h64e6f15e;
    ram_cell[     518] = 32'he30149b6;
    ram_cell[     519] = 32'hcd94ec01;
    ram_cell[     520] = 32'h113f8edc;
    ram_cell[     521] = 32'hf8d4536c;
    ram_cell[     522] = 32'h628b58dc;
    ram_cell[     523] = 32'h9c0b4fb1;
    ram_cell[     524] = 32'h444be981;
    ram_cell[     525] = 32'h4162bc31;
    ram_cell[     526] = 32'hf9c3fcbc;
    ram_cell[     527] = 32'hb7a7c7b9;
    ram_cell[     528] = 32'h369188f9;
    ram_cell[     529] = 32'h1b787604;
    ram_cell[     530] = 32'h004271dc;
    ram_cell[     531] = 32'h6ba40dbf;
    ram_cell[     532] = 32'he4a74005;
    ram_cell[     533] = 32'h95ebe5ba;
    ram_cell[     534] = 32'hdce5b37d;
    ram_cell[     535] = 32'h0794798d;
    ram_cell[     536] = 32'h10dc5a25;
    ram_cell[     537] = 32'hdb2fc150;
    ram_cell[     538] = 32'hf0a59c85;
    ram_cell[     539] = 32'hd6655496;
    ram_cell[     540] = 32'h5a69c440;
    ram_cell[     541] = 32'ha18ea021;
    ram_cell[     542] = 32'h74746109;
    ram_cell[     543] = 32'hf30c0f76;
    ram_cell[     544] = 32'h9408a2c1;
    ram_cell[     545] = 32'h7f534339;
    ram_cell[     546] = 32'he1594f69;
    ram_cell[     547] = 32'h9c378274;
    ram_cell[     548] = 32'h7d991bb5;
    ram_cell[     549] = 32'hc2323578;
    ram_cell[     550] = 32'h81264fd3;
    ram_cell[     551] = 32'hd889751d;
    ram_cell[     552] = 32'hdb30b2c5;
    ram_cell[     553] = 32'he32362ef;
    ram_cell[     554] = 32'hbddc1be5;
    ram_cell[     555] = 32'h59a9e6ac;
    ram_cell[     556] = 32'hf646590e;
    ram_cell[     557] = 32'haf88c554;
    ram_cell[     558] = 32'h13646b14;
    ram_cell[     559] = 32'ha62989d3;
    ram_cell[     560] = 32'h46ae9c07;
    ram_cell[     561] = 32'h4782fc6a;
    ram_cell[     562] = 32'h2d329479;
    ram_cell[     563] = 32'h92f9fa58;
    ram_cell[     564] = 32'hf2a7e694;
    ram_cell[     565] = 32'h74c1cc12;
    ram_cell[     566] = 32'hf795f6f6;
    ram_cell[     567] = 32'h49a88ba2;
    ram_cell[     568] = 32'h63a55fa6;
    ram_cell[     569] = 32'h2904ae6b;
    ram_cell[     570] = 32'hd6878867;
    ram_cell[     571] = 32'hfcbbff41;
    ram_cell[     572] = 32'h2dba60e5;
    ram_cell[     573] = 32'h95bbb079;
    ram_cell[     574] = 32'h51b57fdc;
    ram_cell[     575] = 32'h8d2027bc;
    ram_cell[     576] = 32'hd65aa0c4;
    ram_cell[     577] = 32'h6e0d90ce;
    ram_cell[     578] = 32'h1de1b950;
    ram_cell[     579] = 32'hd9f3ecb9;
    ram_cell[     580] = 32'h70797521;
    ram_cell[     581] = 32'h090cad5a;
    ram_cell[     582] = 32'h77655f9e;
    ram_cell[     583] = 32'h2beb51b2;
    ram_cell[     584] = 32'hefb3adcb;
    ram_cell[     585] = 32'h6072176f;
    ram_cell[     586] = 32'h749819fc;
    ram_cell[     587] = 32'h425a2632;
    ram_cell[     588] = 32'h0e7aecc0;
    ram_cell[     589] = 32'hf1e48ad7;
    ram_cell[     590] = 32'h29e9302d;
    ram_cell[     591] = 32'hf072ed66;
    ram_cell[     592] = 32'hb72ed75a;
    ram_cell[     593] = 32'ha748c708;
    ram_cell[     594] = 32'h1c4e677e;
    ram_cell[     595] = 32'h55fd369f;
    ram_cell[     596] = 32'h5144f7c0;
    ram_cell[     597] = 32'hab52e739;
    ram_cell[     598] = 32'h1820e26f;
    ram_cell[     599] = 32'h214519fb;
    ram_cell[     600] = 32'h53e319df;
    ram_cell[     601] = 32'h66b186b6;
    ram_cell[     602] = 32'hc2dbb80e;
    ram_cell[     603] = 32'h3402a7f0;
    ram_cell[     604] = 32'h4dfe35c7;
    ram_cell[     605] = 32'hc1c4da9a;
    ram_cell[     606] = 32'heb859056;
    ram_cell[     607] = 32'hbfe5e28c;
    ram_cell[     608] = 32'h9d61cc7e;
    ram_cell[     609] = 32'h2666dd20;
    ram_cell[     610] = 32'ha4d741f2;
    ram_cell[     611] = 32'hb1ac83fd;
    ram_cell[     612] = 32'haec1dfe0;
    ram_cell[     613] = 32'h165a7f69;
    ram_cell[     614] = 32'hd1394933;
    ram_cell[     615] = 32'h3039de8e;
    ram_cell[     616] = 32'h50776f26;
    ram_cell[     617] = 32'h8fd06364;
    ram_cell[     618] = 32'hdd9691ae;
    ram_cell[     619] = 32'he2706af8;
    ram_cell[     620] = 32'h56808160;
    ram_cell[     621] = 32'h060471ad;
    ram_cell[     622] = 32'hf38d6835;
    ram_cell[     623] = 32'he8ef741f;
    ram_cell[     624] = 32'h88defff3;
    ram_cell[     625] = 32'h5f6b54d9;
    ram_cell[     626] = 32'h237561d2;
    ram_cell[     627] = 32'h99d7c29b;
    ram_cell[     628] = 32'h2b3e0213;
    ram_cell[     629] = 32'ha257e6de;
    ram_cell[     630] = 32'ha264f956;
    ram_cell[     631] = 32'h47ae9b23;
    ram_cell[     632] = 32'h678c8479;
    ram_cell[     633] = 32'h50deb182;
    ram_cell[     634] = 32'hc8aede93;
    ram_cell[     635] = 32'h971ccc68;
    ram_cell[     636] = 32'h791f4702;
    ram_cell[     637] = 32'h8b1e2fa2;
    ram_cell[     638] = 32'heea0f08d;
    ram_cell[     639] = 32'h03ece7af;
    ram_cell[     640] = 32'hb7f1fc68;
    ram_cell[     641] = 32'hae913ba5;
    ram_cell[     642] = 32'h65e6c180;
    ram_cell[     643] = 32'h62673efc;
    ram_cell[     644] = 32'hb3aa1f18;
    ram_cell[     645] = 32'he728277a;
    ram_cell[     646] = 32'h134c31ee;
    ram_cell[     647] = 32'h17961cae;
    ram_cell[     648] = 32'hf9cbb77b;
    ram_cell[     649] = 32'h5919e1ce;
    ram_cell[     650] = 32'h4ae2ae1e;
    ram_cell[     651] = 32'h5e2be7a4;
    ram_cell[     652] = 32'hb4f94968;
    ram_cell[     653] = 32'h83c6985e;
    ram_cell[     654] = 32'h808be59d;
    ram_cell[     655] = 32'h40032ee2;
    ram_cell[     656] = 32'hb2b595df;
    ram_cell[     657] = 32'h4c63ee0f;
    ram_cell[     658] = 32'hb49f8baa;
    ram_cell[     659] = 32'hde235bc8;
    ram_cell[     660] = 32'h9bbc9fc9;
    ram_cell[     661] = 32'ha72b6d98;
    ram_cell[     662] = 32'h0356ec0b;
    ram_cell[     663] = 32'h4d63a9a0;
    ram_cell[     664] = 32'h2538bec6;
    ram_cell[     665] = 32'h798165ff;
    ram_cell[     666] = 32'h0fa1847d;
    ram_cell[     667] = 32'hd41e6202;
    ram_cell[     668] = 32'h2daf47f7;
    ram_cell[     669] = 32'hac384d2b;
    ram_cell[     670] = 32'h65747cdc;
    ram_cell[     671] = 32'h3ab31c34;
    ram_cell[     672] = 32'h15cf9a6f;
    ram_cell[     673] = 32'he5d98b5b;
    ram_cell[     674] = 32'h3ae47d3c;
    ram_cell[     675] = 32'hfa46e3d6;
    ram_cell[     676] = 32'h03986cf2;
    ram_cell[     677] = 32'h22b74059;
    ram_cell[     678] = 32'hb1d96f50;
    ram_cell[     679] = 32'hfebd0bbf;
    ram_cell[     680] = 32'hd320004e;
    ram_cell[     681] = 32'hd3ed6521;
    ram_cell[     682] = 32'h211be1c2;
    ram_cell[     683] = 32'h9e512e54;
    ram_cell[     684] = 32'hcc3b605e;
    ram_cell[     685] = 32'hf8667be7;
    ram_cell[     686] = 32'h0944c7f7;
    ram_cell[     687] = 32'h4c49b758;
    ram_cell[     688] = 32'haf786ee4;
    ram_cell[     689] = 32'he0c2bf10;
    ram_cell[     690] = 32'h06588919;
    ram_cell[     691] = 32'h366faa33;
    ram_cell[     692] = 32'h983f8529;
    ram_cell[     693] = 32'h5aa949f8;
    ram_cell[     694] = 32'h6bbf28c5;
    ram_cell[     695] = 32'h9ab6c70c;
    ram_cell[     696] = 32'h7839e2d8;
    ram_cell[     697] = 32'h17f2be44;
    ram_cell[     698] = 32'h667b1f88;
    ram_cell[     699] = 32'hd8b07178;
    ram_cell[     700] = 32'h0aba595e;
    ram_cell[     701] = 32'h7fd61445;
    ram_cell[     702] = 32'h92bf5a69;
    ram_cell[     703] = 32'hd4fa2354;
    ram_cell[     704] = 32'h25102879;
    ram_cell[     705] = 32'h7f7a83c4;
    ram_cell[     706] = 32'h078c44c4;
    ram_cell[     707] = 32'h77bc7347;
    ram_cell[     708] = 32'h11e392bd;
    ram_cell[     709] = 32'heff8e9d1;
    ram_cell[     710] = 32'h62240988;
    ram_cell[     711] = 32'h7ec37d10;
    ram_cell[     712] = 32'h75a02eac;
    ram_cell[     713] = 32'h76989168;
    ram_cell[     714] = 32'h4727e362;
    ram_cell[     715] = 32'h94e50cb2;
    ram_cell[     716] = 32'he0a88525;
    ram_cell[     717] = 32'hf12c1506;
    ram_cell[     718] = 32'h71d2dcf3;
    ram_cell[     719] = 32'h71cc7278;
    ram_cell[     720] = 32'h657b4843;
    ram_cell[     721] = 32'h70d2443c;
    ram_cell[     722] = 32'h9a37af73;
    ram_cell[     723] = 32'hd97b924d;
    ram_cell[     724] = 32'h2bdccc44;
    ram_cell[     725] = 32'hea9887d6;
    ram_cell[     726] = 32'h15fb0580;
    ram_cell[     727] = 32'h7d00208d;
    ram_cell[     728] = 32'he07ada7e;
    ram_cell[     729] = 32'h7306383a;
    ram_cell[     730] = 32'h961767d5;
    ram_cell[     731] = 32'hf8f79b69;
    ram_cell[     732] = 32'hfda733ca;
    ram_cell[     733] = 32'hf8691414;
    ram_cell[     734] = 32'heccf8c66;
    ram_cell[     735] = 32'h192b362b;
    ram_cell[     736] = 32'hd87fe8d3;
    ram_cell[     737] = 32'hd40b76ad;
    ram_cell[     738] = 32'he16b2629;
    ram_cell[     739] = 32'hb45a55a8;
    ram_cell[     740] = 32'hdeb65e65;
    ram_cell[     741] = 32'h261d8c04;
    ram_cell[     742] = 32'haa6cd7da;
    ram_cell[     743] = 32'h4694c0dd;
    ram_cell[     744] = 32'hf391d8c9;
    ram_cell[     745] = 32'h54459296;
    ram_cell[     746] = 32'h0fe978a3;
    ram_cell[     747] = 32'h3e883dfa;
    ram_cell[     748] = 32'hbd41bbcf;
    ram_cell[     749] = 32'h0b47e802;
    ram_cell[     750] = 32'hef388ac3;
    ram_cell[     751] = 32'h2cf403a9;
    ram_cell[     752] = 32'h696150ed;
    ram_cell[     753] = 32'h986415cd;
    ram_cell[     754] = 32'h536cfd6b;
    ram_cell[     755] = 32'h7b21a968;
    ram_cell[     756] = 32'h0a7007b9;
    ram_cell[     757] = 32'h42e89020;
    ram_cell[     758] = 32'h0082e76d;
    ram_cell[     759] = 32'h85414eec;
    ram_cell[     760] = 32'h92296fb2;
    ram_cell[     761] = 32'h8f82f04b;
    ram_cell[     762] = 32'h7177474e;
    ram_cell[     763] = 32'h8418dae9;
    ram_cell[     764] = 32'h4bf67d43;
    ram_cell[     765] = 32'hf76b6e8e;
    ram_cell[     766] = 32'h9c756e45;
    ram_cell[     767] = 32'ha2e2c726;
end

endmodule

