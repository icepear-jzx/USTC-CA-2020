
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h797743d7;
    ram_cell[       1] = 32'h0;  // 32'h36b89901;
    ram_cell[       2] = 32'h0;  // 32'h035fdc9a;
    ram_cell[       3] = 32'h0;  // 32'ha28c0f99;
    ram_cell[       4] = 32'h0;  // 32'h08d8cded;
    ram_cell[       5] = 32'h0;  // 32'h1a10afac;
    ram_cell[       6] = 32'h0;  // 32'h7359c785;
    ram_cell[       7] = 32'h0;  // 32'ha11bb49d;
    ram_cell[       8] = 32'h0;  // 32'h9b9a4db7;
    ram_cell[       9] = 32'h0;  // 32'ha427b5f6;
    ram_cell[      10] = 32'h0;  // 32'h44847363;
    ram_cell[      11] = 32'h0;  // 32'h98f767ed;
    ram_cell[      12] = 32'h0;  // 32'h1694ce3d;
    ram_cell[      13] = 32'h0;  // 32'h26365b7b;
    ram_cell[      14] = 32'h0;  // 32'h2007093c;
    ram_cell[      15] = 32'h0;  // 32'h19e8e946;
    ram_cell[      16] = 32'h0;  // 32'hb9a0d76b;
    ram_cell[      17] = 32'h0;  // 32'h8483c94b;
    ram_cell[      18] = 32'h0;  // 32'hb68d5699;
    ram_cell[      19] = 32'h0;  // 32'h14d2c6b9;
    ram_cell[      20] = 32'h0;  // 32'hc97a4b6b;
    ram_cell[      21] = 32'h0;  // 32'h43211874;
    ram_cell[      22] = 32'h0;  // 32'hb9ad3d36;
    ram_cell[      23] = 32'h0;  // 32'hfbfa06b9;
    ram_cell[      24] = 32'h0;  // 32'hbfbe0546;
    ram_cell[      25] = 32'h0;  // 32'h2373b879;
    ram_cell[      26] = 32'h0;  // 32'he3885c27;
    ram_cell[      27] = 32'h0;  // 32'hffe3436d;
    ram_cell[      28] = 32'h0;  // 32'h25d2a7ec;
    ram_cell[      29] = 32'h0;  // 32'h965f31d0;
    ram_cell[      30] = 32'h0;  // 32'h4f2533f1;
    ram_cell[      31] = 32'h0;  // 32'ha17f98d4;
    ram_cell[      32] = 32'h0;  // 32'h4c5ff3bd;
    ram_cell[      33] = 32'h0;  // 32'h58f4f321;
    ram_cell[      34] = 32'h0;  // 32'h35d08f8c;
    ram_cell[      35] = 32'h0;  // 32'hecfb2880;
    ram_cell[      36] = 32'h0;  // 32'h2184568f;
    ram_cell[      37] = 32'h0;  // 32'h02bdf270;
    ram_cell[      38] = 32'h0;  // 32'h7a9790b4;
    ram_cell[      39] = 32'h0;  // 32'h0a073238;
    ram_cell[      40] = 32'h0;  // 32'h48e14737;
    ram_cell[      41] = 32'h0;  // 32'hf9b627ce;
    ram_cell[      42] = 32'h0;  // 32'h01b131c6;
    ram_cell[      43] = 32'h0;  // 32'hf2307b53;
    ram_cell[      44] = 32'h0;  // 32'he775d4fa;
    ram_cell[      45] = 32'h0;  // 32'he7496da9;
    ram_cell[      46] = 32'h0;  // 32'ha998073e;
    ram_cell[      47] = 32'h0;  // 32'h86d658c2;
    ram_cell[      48] = 32'h0;  // 32'h9e0887c6;
    ram_cell[      49] = 32'h0;  // 32'h8e69a03c;
    ram_cell[      50] = 32'h0;  // 32'hc0331622;
    ram_cell[      51] = 32'h0;  // 32'hc569fb14;
    ram_cell[      52] = 32'h0;  // 32'hfb1a3698;
    ram_cell[      53] = 32'h0;  // 32'hd00fb76d;
    ram_cell[      54] = 32'h0;  // 32'heec8e519;
    ram_cell[      55] = 32'h0;  // 32'h63b09f93;
    ram_cell[      56] = 32'h0;  // 32'hd9d87b38;
    ram_cell[      57] = 32'h0;  // 32'hdacd98dd;
    ram_cell[      58] = 32'h0;  // 32'hf1f9662b;
    ram_cell[      59] = 32'h0;  // 32'h77d9202d;
    ram_cell[      60] = 32'h0;  // 32'he4de9bdd;
    ram_cell[      61] = 32'h0;  // 32'h867176d4;
    ram_cell[      62] = 32'h0;  // 32'h64021d30;
    ram_cell[      63] = 32'h0;  // 32'h49d1649e;
    ram_cell[      64] = 32'h0;  // 32'h6e7359cf;
    ram_cell[      65] = 32'h0;  // 32'h3d81c82f;
    ram_cell[      66] = 32'h0;  // 32'h5f2065d9;
    ram_cell[      67] = 32'h0;  // 32'h514a5236;
    ram_cell[      68] = 32'h0;  // 32'h8608437e;
    ram_cell[      69] = 32'h0;  // 32'he4a14800;
    ram_cell[      70] = 32'h0;  // 32'h5ccb71f4;
    ram_cell[      71] = 32'h0;  // 32'h694fbc7a;
    ram_cell[      72] = 32'h0;  // 32'h8e3d566c;
    ram_cell[      73] = 32'h0;  // 32'h52359498;
    ram_cell[      74] = 32'h0;  // 32'h8109f364;
    ram_cell[      75] = 32'h0;  // 32'hea0c4150;
    ram_cell[      76] = 32'h0;  // 32'h172f46ca;
    ram_cell[      77] = 32'h0;  // 32'h34ba003c;
    ram_cell[      78] = 32'h0;  // 32'h0f94c278;
    ram_cell[      79] = 32'h0;  // 32'h3617e34b;
    ram_cell[      80] = 32'h0;  // 32'h68ac6b9e;
    ram_cell[      81] = 32'h0;  // 32'h40436f14;
    ram_cell[      82] = 32'h0;  // 32'h20bd2849;
    ram_cell[      83] = 32'h0;  // 32'h4b129eb7;
    ram_cell[      84] = 32'h0;  // 32'ha69f31de;
    ram_cell[      85] = 32'h0;  // 32'h0c8eac84;
    ram_cell[      86] = 32'h0;  // 32'he69ecd31;
    ram_cell[      87] = 32'h0;  // 32'h129368d3;
    ram_cell[      88] = 32'h0;  // 32'h9eb9931c;
    ram_cell[      89] = 32'h0;  // 32'hc9d8bf75;
    ram_cell[      90] = 32'h0;  // 32'h6e173cd0;
    ram_cell[      91] = 32'h0;  // 32'h66988ad8;
    ram_cell[      92] = 32'h0;  // 32'hdedba05d;
    ram_cell[      93] = 32'h0;  // 32'h17e47e9b;
    ram_cell[      94] = 32'h0;  // 32'hb3998a97;
    ram_cell[      95] = 32'h0;  // 32'h5ff25765;
    ram_cell[      96] = 32'h0;  // 32'h66c70ecf;
    ram_cell[      97] = 32'h0;  // 32'hef7c1bca;
    ram_cell[      98] = 32'h0;  // 32'hf1235b4e;
    ram_cell[      99] = 32'h0;  // 32'hb0e88c84;
    ram_cell[     100] = 32'h0;  // 32'hee9dc659;
    ram_cell[     101] = 32'h0;  // 32'h9dd34fa4;
    ram_cell[     102] = 32'h0;  // 32'hcaaf6e30;
    ram_cell[     103] = 32'h0;  // 32'h0004a43b;
    ram_cell[     104] = 32'h0;  // 32'heca9cca8;
    ram_cell[     105] = 32'h0;  // 32'ha64f8cd7;
    ram_cell[     106] = 32'h0;  // 32'h2e143334;
    ram_cell[     107] = 32'h0;  // 32'h1ccaeb8f;
    ram_cell[     108] = 32'h0;  // 32'h828762c2;
    ram_cell[     109] = 32'h0;  // 32'h57ad05b2;
    ram_cell[     110] = 32'h0;  // 32'hb67e99ad;
    ram_cell[     111] = 32'h0;  // 32'h9fe8e500;
    ram_cell[     112] = 32'h0;  // 32'h15c100d2;
    ram_cell[     113] = 32'h0;  // 32'hb4444c06;
    ram_cell[     114] = 32'h0;  // 32'hedd72c86;
    ram_cell[     115] = 32'h0;  // 32'h6a8fd15d;
    ram_cell[     116] = 32'h0;  // 32'ha435f044;
    ram_cell[     117] = 32'h0;  // 32'hb8df2346;
    ram_cell[     118] = 32'h0;  // 32'h9a615ee4;
    ram_cell[     119] = 32'h0;  // 32'h8fe689fb;
    ram_cell[     120] = 32'h0;  // 32'h0a3f9edf;
    ram_cell[     121] = 32'h0;  // 32'h760b0dce;
    ram_cell[     122] = 32'h0;  // 32'hfc5bedc2;
    ram_cell[     123] = 32'h0;  // 32'had10b1e0;
    ram_cell[     124] = 32'h0;  // 32'h872adffe;
    ram_cell[     125] = 32'h0;  // 32'hf72a97a7;
    ram_cell[     126] = 32'h0;  // 32'h6e84cf1a;
    ram_cell[     127] = 32'h0;  // 32'h43a23d8b;
    ram_cell[     128] = 32'h0;  // 32'h715fea76;
    ram_cell[     129] = 32'h0;  // 32'h12ed1607;
    ram_cell[     130] = 32'h0;  // 32'h54394ad9;
    ram_cell[     131] = 32'h0;  // 32'h3cb6d9cc;
    ram_cell[     132] = 32'h0;  // 32'h6e35574f;
    ram_cell[     133] = 32'h0;  // 32'hd2e9621e;
    ram_cell[     134] = 32'h0;  // 32'h6445baf9;
    ram_cell[     135] = 32'h0;  // 32'h4c881d3d;
    ram_cell[     136] = 32'h0;  // 32'hbec0eefa;
    ram_cell[     137] = 32'h0;  // 32'h7ca9d032;
    ram_cell[     138] = 32'h0;  // 32'hc8967006;
    ram_cell[     139] = 32'h0;  // 32'h38c47cdc;
    ram_cell[     140] = 32'h0;  // 32'hbbb7e568;
    ram_cell[     141] = 32'h0;  // 32'he4ad7953;
    ram_cell[     142] = 32'h0;  // 32'h07dd47dd;
    ram_cell[     143] = 32'h0;  // 32'hd147ba90;
    ram_cell[     144] = 32'h0;  // 32'hb12cfbe8;
    ram_cell[     145] = 32'h0;  // 32'h79e6939e;
    ram_cell[     146] = 32'h0;  // 32'hc02629b5;
    ram_cell[     147] = 32'h0;  // 32'h6af87a84;
    ram_cell[     148] = 32'h0;  // 32'h0dc1dffc;
    ram_cell[     149] = 32'h0;  // 32'h8841de1a;
    ram_cell[     150] = 32'h0;  // 32'h646155fe;
    ram_cell[     151] = 32'h0;  // 32'h010507db;
    ram_cell[     152] = 32'h0;  // 32'hdbb805ac;
    ram_cell[     153] = 32'h0;  // 32'h98a16341;
    ram_cell[     154] = 32'h0;  // 32'h7b5b218e;
    ram_cell[     155] = 32'h0;  // 32'h1f91d727;
    ram_cell[     156] = 32'h0;  // 32'he73616d8;
    ram_cell[     157] = 32'h0;  // 32'hed5db0fd;
    ram_cell[     158] = 32'h0;  // 32'h910bcc6c;
    ram_cell[     159] = 32'h0;  // 32'hc504706a;
    ram_cell[     160] = 32'h0;  // 32'hb88823c2;
    ram_cell[     161] = 32'h0;  // 32'ha80e5206;
    ram_cell[     162] = 32'h0;  // 32'ha14717cd;
    ram_cell[     163] = 32'h0;  // 32'h80138547;
    ram_cell[     164] = 32'h0;  // 32'h96a167b2;
    ram_cell[     165] = 32'h0;  // 32'ha28951f2;
    ram_cell[     166] = 32'h0;  // 32'h0b5f31b4;
    ram_cell[     167] = 32'h0;  // 32'h305aab3e;
    ram_cell[     168] = 32'h0;  // 32'h721f6364;
    ram_cell[     169] = 32'h0;  // 32'hcede20c5;
    ram_cell[     170] = 32'h0;  // 32'h76e26987;
    ram_cell[     171] = 32'h0;  // 32'hd75e7d0d;
    ram_cell[     172] = 32'h0;  // 32'h8c46dba1;
    ram_cell[     173] = 32'h0;  // 32'haee6b371;
    ram_cell[     174] = 32'h0;  // 32'h9904e6e5;
    ram_cell[     175] = 32'h0;  // 32'hb0df9ab5;
    ram_cell[     176] = 32'h0;  // 32'hea7e6231;
    ram_cell[     177] = 32'h0;  // 32'hfba1746d;
    ram_cell[     178] = 32'h0;  // 32'h002e04e1;
    ram_cell[     179] = 32'h0;  // 32'hd166e0ba;
    ram_cell[     180] = 32'h0;  // 32'h24bf3c3f;
    ram_cell[     181] = 32'h0;  // 32'h3270dcec;
    ram_cell[     182] = 32'h0;  // 32'hbc853ebf;
    ram_cell[     183] = 32'h0;  // 32'hdac850f0;
    ram_cell[     184] = 32'h0;  // 32'h0e6a87ce;
    ram_cell[     185] = 32'h0;  // 32'h381c0872;
    ram_cell[     186] = 32'h0;  // 32'h58182599;
    ram_cell[     187] = 32'h0;  // 32'h921a2770;
    ram_cell[     188] = 32'h0;  // 32'hd909c204;
    ram_cell[     189] = 32'h0;  // 32'h0eb14f2d;
    ram_cell[     190] = 32'h0;  // 32'h0b719805;
    ram_cell[     191] = 32'h0;  // 32'h851e64da;
    ram_cell[     192] = 32'h0;  // 32'h12e9ce7d;
    ram_cell[     193] = 32'h0;  // 32'he2061e27;
    ram_cell[     194] = 32'h0;  // 32'hb2fb85b2;
    ram_cell[     195] = 32'h0;  // 32'hbcd48651;
    ram_cell[     196] = 32'h0;  // 32'h42e0315c;
    ram_cell[     197] = 32'h0;  // 32'h96cc6a77;
    ram_cell[     198] = 32'h0;  // 32'h64be958d;
    ram_cell[     199] = 32'h0;  // 32'h8d61b1e8;
    ram_cell[     200] = 32'h0;  // 32'h09ec40df;
    ram_cell[     201] = 32'h0;  // 32'h4ad0cff9;
    ram_cell[     202] = 32'h0;  // 32'hc5355576;
    ram_cell[     203] = 32'h0;  // 32'h73366b6b;
    ram_cell[     204] = 32'h0;  // 32'hfe8a6946;
    ram_cell[     205] = 32'h0;  // 32'hef871151;
    ram_cell[     206] = 32'h0;  // 32'h4a327142;
    ram_cell[     207] = 32'h0;  // 32'h3aabef6f;
    ram_cell[     208] = 32'h0;  // 32'h1477ef18;
    ram_cell[     209] = 32'h0;  // 32'h79d5525f;
    ram_cell[     210] = 32'h0;  // 32'h427b01d2;
    ram_cell[     211] = 32'h0;  // 32'h4f06b9f1;
    ram_cell[     212] = 32'h0;  // 32'h4b76b7a1;
    ram_cell[     213] = 32'h0;  // 32'ha36b38f7;
    ram_cell[     214] = 32'h0;  // 32'h53b146ef;
    ram_cell[     215] = 32'h0;  // 32'h9d434527;
    ram_cell[     216] = 32'h0;  // 32'h9d274182;
    ram_cell[     217] = 32'h0;  // 32'hac812e9f;
    ram_cell[     218] = 32'h0;  // 32'h0239e3af;
    ram_cell[     219] = 32'h0;  // 32'h49b9bbd2;
    ram_cell[     220] = 32'h0;  // 32'h2e576ec3;
    ram_cell[     221] = 32'h0;  // 32'h13f4c775;
    ram_cell[     222] = 32'h0;  // 32'h295ac5ca;
    ram_cell[     223] = 32'h0;  // 32'ha2117b9d;
    ram_cell[     224] = 32'h0;  // 32'h34ba771e;
    ram_cell[     225] = 32'h0;  // 32'h26e7f357;
    ram_cell[     226] = 32'h0;  // 32'he6e0560b;
    ram_cell[     227] = 32'h0;  // 32'he1bac6cc;
    ram_cell[     228] = 32'h0;  // 32'hfb4b1223;
    ram_cell[     229] = 32'h0;  // 32'hbeae9845;
    ram_cell[     230] = 32'h0;  // 32'h7835d440;
    ram_cell[     231] = 32'h0;  // 32'hfe10ea47;
    ram_cell[     232] = 32'h0;  // 32'haa8608ab;
    ram_cell[     233] = 32'h0;  // 32'h6b8312b0;
    ram_cell[     234] = 32'h0;  // 32'heacd485a;
    ram_cell[     235] = 32'h0;  // 32'h33ddcd8c;
    ram_cell[     236] = 32'h0;  // 32'h91c22142;
    ram_cell[     237] = 32'h0;  // 32'ha6445568;
    ram_cell[     238] = 32'h0;  // 32'ha244c53b;
    ram_cell[     239] = 32'h0;  // 32'hfff6ae71;
    ram_cell[     240] = 32'h0;  // 32'h61b4714e;
    ram_cell[     241] = 32'h0;  // 32'hb61ff5c0;
    ram_cell[     242] = 32'h0;  // 32'h88550226;
    ram_cell[     243] = 32'h0;  // 32'h5ee5ecb7;
    ram_cell[     244] = 32'h0;  // 32'h44a75e83;
    ram_cell[     245] = 32'h0;  // 32'h79baf947;
    ram_cell[     246] = 32'h0;  // 32'hfd157a27;
    ram_cell[     247] = 32'h0;  // 32'h59072fba;
    ram_cell[     248] = 32'h0;  // 32'hb1a8ff62;
    ram_cell[     249] = 32'h0;  // 32'hf4e92bd0;
    ram_cell[     250] = 32'h0;  // 32'he4041a50;
    ram_cell[     251] = 32'h0;  // 32'h3959e283;
    ram_cell[     252] = 32'h0;  // 32'h7d42c394;
    ram_cell[     253] = 32'h0;  // 32'h04b0557f;
    ram_cell[     254] = 32'h0;  // 32'h58f68363;
    ram_cell[     255] = 32'h0;  // 32'h0a2c8678;
    ram_cell[     256] = 32'h0;  // 32'h2281d20f;
    ram_cell[     257] = 32'h0;  // 32'h4630da2c;
    ram_cell[     258] = 32'h0;  // 32'he38b7db2;
    ram_cell[     259] = 32'h0;  // 32'h1e293588;
    ram_cell[     260] = 32'h0;  // 32'h761eb690;
    ram_cell[     261] = 32'h0;  // 32'h9a3cbbed;
    ram_cell[     262] = 32'h0;  // 32'h7e8d005e;
    ram_cell[     263] = 32'h0;  // 32'h3693c4bf;
    ram_cell[     264] = 32'h0;  // 32'hb4450560;
    ram_cell[     265] = 32'h0;  // 32'h9361e8df;
    ram_cell[     266] = 32'h0;  // 32'hfcd1f44f;
    ram_cell[     267] = 32'h0;  // 32'h5a34756a;
    ram_cell[     268] = 32'h0;  // 32'h63126af2;
    ram_cell[     269] = 32'h0;  // 32'hfc16b295;
    ram_cell[     270] = 32'h0;  // 32'hbdfa1587;
    ram_cell[     271] = 32'h0;  // 32'h9b48d742;
    ram_cell[     272] = 32'h0;  // 32'h43c421c4;
    ram_cell[     273] = 32'h0;  // 32'haddd6478;
    ram_cell[     274] = 32'h0;  // 32'hcd0a664c;
    ram_cell[     275] = 32'h0;  // 32'h4d9d894c;
    ram_cell[     276] = 32'h0;  // 32'h43905b35;
    ram_cell[     277] = 32'h0;  // 32'hc70e9897;
    ram_cell[     278] = 32'h0;  // 32'he630fb89;
    ram_cell[     279] = 32'h0;  // 32'hfeb52db8;
    ram_cell[     280] = 32'h0;  // 32'hbd7347f2;
    ram_cell[     281] = 32'h0;  // 32'hf53d71c9;
    ram_cell[     282] = 32'h0;  // 32'h2b9dad31;
    ram_cell[     283] = 32'h0;  // 32'h29ae26a1;
    ram_cell[     284] = 32'h0;  // 32'h8ac08f62;
    ram_cell[     285] = 32'h0;  // 32'hca41b586;
    ram_cell[     286] = 32'h0;  // 32'h209d046f;
    ram_cell[     287] = 32'h0;  // 32'haa417aa8;
    ram_cell[     288] = 32'h0;  // 32'hc54c753c;
    ram_cell[     289] = 32'h0;  // 32'h6f9ba051;
    ram_cell[     290] = 32'h0;  // 32'h94fbab6d;
    ram_cell[     291] = 32'h0;  // 32'hb4afbd39;
    ram_cell[     292] = 32'h0;  // 32'hbf8b7c01;
    ram_cell[     293] = 32'h0;  // 32'h74924951;
    ram_cell[     294] = 32'h0;  // 32'h0d563749;
    ram_cell[     295] = 32'h0;  // 32'hb8ff1b26;
    ram_cell[     296] = 32'h0;  // 32'h3101cb58;
    ram_cell[     297] = 32'h0;  // 32'ha63da01a;
    ram_cell[     298] = 32'h0;  // 32'hc8a6c80f;
    ram_cell[     299] = 32'h0;  // 32'hb2536f69;
    ram_cell[     300] = 32'h0;  // 32'h75d0ab5c;
    ram_cell[     301] = 32'h0;  // 32'h2d824079;
    ram_cell[     302] = 32'h0;  // 32'hf46b1358;
    ram_cell[     303] = 32'h0;  // 32'h673555e5;
    ram_cell[     304] = 32'h0;  // 32'h3da7290e;
    ram_cell[     305] = 32'h0;  // 32'h0a302d97;
    ram_cell[     306] = 32'h0;  // 32'hbbbee080;
    ram_cell[     307] = 32'h0;  // 32'h0802cf37;
    ram_cell[     308] = 32'h0;  // 32'ha480b199;
    ram_cell[     309] = 32'h0;  // 32'he7bf7dfb;
    ram_cell[     310] = 32'h0;  // 32'h6f7d40c0;
    ram_cell[     311] = 32'h0;  // 32'hb909becb;
    ram_cell[     312] = 32'h0;  // 32'h77409799;
    ram_cell[     313] = 32'h0;  // 32'h9f73a89a;
    ram_cell[     314] = 32'h0;  // 32'h1732acb6;
    ram_cell[     315] = 32'h0;  // 32'h1bed2df8;
    ram_cell[     316] = 32'h0;  // 32'h55cb033b;
    ram_cell[     317] = 32'h0;  // 32'h5c55396c;
    ram_cell[     318] = 32'h0;  // 32'hbdb31047;
    ram_cell[     319] = 32'h0;  // 32'hb3aecee7;
    ram_cell[     320] = 32'h0;  // 32'h54705086;
    ram_cell[     321] = 32'h0;  // 32'h22b2d612;
    ram_cell[     322] = 32'h0;  // 32'h61b591bb;
    ram_cell[     323] = 32'h0;  // 32'hcb94ae6e;
    ram_cell[     324] = 32'h0;  // 32'h3960d35c;
    ram_cell[     325] = 32'h0;  // 32'h52c8da13;
    ram_cell[     326] = 32'h0;  // 32'h8650c7cb;
    ram_cell[     327] = 32'h0;  // 32'he8431e08;
    ram_cell[     328] = 32'h0;  // 32'h6c1ded89;
    ram_cell[     329] = 32'h0;  // 32'hec076454;
    ram_cell[     330] = 32'h0;  // 32'h5821a96e;
    ram_cell[     331] = 32'h0;  // 32'h3efeb05c;
    ram_cell[     332] = 32'h0;  // 32'hade2f1ae;
    ram_cell[     333] = 32'h0;  // 32'h2f0389bf;
    ram_cell[     334] = 32'h0;  // 32'h72740fed;
    ram_cell[     335] = 32'h0;  // 32'he029282d;
    ram_cell[     336] = 32'h0;  // 32'h15ccc5df;
    ram_cell[     337] = 32'h0;  // 32'h98a627d0;
    ram_cell[     338] = 32'h0;  // 32'h398c6a47;
    ram_cell[     339] = 32'h0;  // 32'h220749e4;
    ram_cell[     340] = 32'h0;  // 32'h135529bf;
    ram_cell[     341] = 32'h0;  // 32'h523b24da;
    ram_cell[     342] = 32'h0;  // 32'h69b3397e;
    ram_cell[     343] = 32'h0;  // 32'hf66298c3;
    ram_cell[     344] = 32'h0;  // 32'h050fc9ef;
    ram_cell[     345] = 32'h0;  // 32'h044ffb31;
    ram_cell[     346] = 32'h0;  // 32'h8cb08437;
    ram_cell[     347] = 32'h0;  // 32'h4d3204e2;
    ram_cell[     348] = 32'h0;  // 32'h0f77bf6f;
    ram_cell[     349] = 32'h0;  // 32'h11513415;
    ram_cell[     350] = 32'h0;  // 32'he597c511;
    ram_cell[     351] = 32'h0;  // 32'h5e521393;
    ram_cell[     352] = 32'h0;  // 32'h8a6f5327;
    ram_cell[     353] = 32'h0;  // 32'h0befa29c;
    ram_cell[     354] = 32'h0;  // 32'ha88b11da;
    ram_cell[     355] = 32'h0;  // 32'h6af9856f;
    ram_cell[     356] = 32'h0;  // 32'h7d46c0ad;
    ram_cell[     357] = 32'h0;  // 32'hc12cf38f;
    ram_cell[     358] = 32'h0;  // 32'hedf28435;
    ram_cell[     359] = 32'h0;  // 32'h58003d82;
    ram_cell[     360] = 32'h0;  // 32'h51c74930;
    ram_cell[     361] = 32'h0;  // 32'h5e60d32e;
    ram_cell[     362] = 32'h0;  // 32'hc1083ba0;
    ram_cell[     363] = 32'h0;  // 32'hec5b47f7;
    ram_cell[     364] = 32'h0;  // 32'h7a1bfe67;
    ram_cell[     365] = 32'h0;  // 32'h2e1a2a3f;
    ram_cell[     366] = 32'h0;  // 32'h7b0e5ac9;
    ram_cell[     367] = 32'h0;  // 32'h30ace3f2;
    ram_cell[     368] = 32'h0;  // 32'ha4a14291;
    ram_cell[     369] = 32'h0;  // 32'hbe6c382f;
    ram_cell[     370] = 32'h0;  // 32'h21b3926a;
    ram_cell[     371] = 32'h0;  // 32'h6b5473c2;
    ram_cell[     372] = 32'h0;  // 32'hf4e0b97d;
    ram_cell[     373] = 32'h0;  // 32'h9d38bd88;
    ram_cell[     374] = 32'h0;  // 32'hea82dcb6;
    ram_cell[     375] = 32'h0;  // 32'hb908b431;
    ram_cell[     376] = 32'h0;  // 32'hb6176d31;
    ram_cell[     377] = 32'h0;  // 32'h29ff83d3;
    ram_cell[     378] = 32'h0;  // 32'hba6c2532;
    ram_cell[     379] = 32'h0;  // 32'hd420f038;
    ram_cell[     380] = 32'h0;  // 32'hf56c8218;
    ram_cell[     381] = 32'h0;  // 32'h7d725197;
    ram_cell[     382] = 32'h0;  // 32'h3942eadb;
    ram_cell[     383] = 32'h0;  // 32'h547efb6f;
    ram_cell[     384] = 32'h0;  // 32'heaca72d8;
    ram_cell[     385] = 32'h0;  // 32'h711b0594;
    ram_cell[     386] = 32'h0;  // 32'h5d132fff;
    ram_cell[     387] = 32'h0;  // 32'h0a5f53e4;
    ram_cell[     388] = 32'h0;  // 32'h1bc6c718;
    ram_cell[     389] = 32'h0;  // 32'h3dd1572d;
    ram_cell[     390] = 32'h0;  // 32'h2cebe520;
    ram_cell[     391] = 32'h0;  // 32'haf480304;
    ram_cell[     392] = 32'h0;  // 32'h0d9addf8;
    ram_cell[     393] = 32'h0;  // 32'h7957f708;
    ram_cell[     394] = 32'h0;  // 32'h0417b8d2;
    ram_cell[     395] = 32'h0;  // 32'h8c315db7;
    ram_cell[     396] = 32'h0;  // 32'hb94777d0;
    ram_cell[     397] = 32'h0;  // 32'ha64731b9;
    ram_cell[     398] = 32'h0;  // 32'h4df69a41;
    ram_cell[     399] = 32'h0;  // 32'h7b6d9745;
    ram_cell[     400] = 32'h0;  // 32'h9d639050;
    ram_cell[     401] = 32'h0;  // 32'h45416d0b;
    ram_cell[     402] = 32'h0;  // 32'h2363e2b6;
    ram_cell[     403] = 32'h0;  // 32'h7bb20913;
    ram_cell[     404] = 32'h0;  // 32'hcd814026;
    ram_cell[     405] = 32'h0;  // 32'habe9b101;
    ram_cell[     406] = 32'h0;  // 32'hb272be3f;
    ram_cell[     407] = 32'h0;  // 32'h63626c16;
    ram_cell[     408] = 32'h0;  // 32'h8cc8796b;
    ram_cell[     409] = 32'h0;  // 32'h836002b0;
    ram_cell[     410] = 32'h0;  // 32'hefee2d48;
    ram_cell[     411] = 32'h0;  // 32'haaf7be3b;
    ram_cell[     412] = 32'h0;  // 32'h4473d12e;
    ram_cell[     413] = 32'h0;  // 32'hc3a79bec;
    ram_cell[     414] = 32'h0;  // 32'h3224b539;
    ram_cell[     415] = 32'h0;  // 32'h2faf52ff;
    ram_cell[     416] = 32'h0;  // 32'he11130c0;
    ram_cell[     417] = 32'h0;  // 32'h954a4f8a;
    ram_cell[     418] = 32'h0;  // 32'h17f35a05;
    ram_cell[     419] = 32'h0;  // 32'h2deb901a;
    ram_cell[     420] = 32'h0;  // 32'h000ebe47;
    ram_cell[     421] = 32'h0;  // 32'h28008742;
    ram_cell[     422] = 32'h0;  // 32'h65817be6;
    ram_cell[     423] = 32'h0;  // 32'hd5dede51;
    ram_cell[     424] = 32'h0;  // 32'h95d74ffa;
    ram_cell[     425] = 32'h0;  // 32'h2ce8ecac;
    ram_cell[     426] = 32'h0;  // 32'h1c80ceb5;
    ram_cell[     427] = 32'h0;  // 32'hf2ec358e;
    ram_cell[     428] = 32'h0;  // 32'h0adc4cc2;
    ram_cell[     429] = 32'h0;  // 32'h9039bce3;
    ram_cell[     430] = 32'h0;  // 32'hafcbf19f;
    ram_cell[     431] = 32'h0;  // 32'he31d922a;
    ram_cell[     432] = 32'h0;  // 32'he299f4dd;
    ram_cell[     433] = 32'h0;  // 32'h531763d7;
    ram_cell[     434] = 32'h0;  // 32'hf21cd4bd;
    ram_cell[     435] = 32'h0;  // 32'hb6f2f90e;
    ram_cell[     436] = 32'h0;  // 32'he53541bf;
    ram_cell[     437] = 32'h0;  // 32'h091afa06;
    ram_cell[     438] = 32'h0;  // 32'h017d105f;
    ram_cell[     439] = 32'h0;  // 32'hf7378f53;
    ram_cell[     440] = 32'h0;  // 32'h2b2bfafa;
    ram_cell[     441] = 32'h0;  // 32'hd3769897;
    ram_cell[     442] = 32'h0;  // 32'h23639512;
    ram_cell[     443] = 32'h0;  // 32'h958b0c0f;
    ram_cell[     444] = 32'h0;  // 32'hb4d2404b;
    ram_cell[     445] = 32'h0;  // 32'hdfed5fc9;
    ram_cell[     446] = 32'h0;  // 32'h3d907fb1;
    ram_cell[     447] = 32'h0;  // 32'hdc97eb9d;
    ram_cell[     448] = 32'h0;  // 32'h9cb38cbc;
    ram_cell[     449] = 32'h0;  // 32'h6e9faa2d;
    ram_cell[     450] = 32'h0;  // 32'h07fba0ae;
    ram_cell[     451] = 32'h0;  // 32'had031ba5;
    ram_cell[     452] = 32'h0;  // 32'hbd04269f;
    ram_cell[     453] = 32'h0;  // 32'h67d179e7;
    ram_cell[     454] = 32'h0;  // 32'h3c0b6239;
    ram_cell[     455] = 32'h0;  // 32'h321a6aa0;
    ram_cell[     456] = 32'h0;  // 32'he417fad2;
    ram_cell[     457] = 32'h0;  // 32'h10ad5651;
    ram_cell[     458] = 32'h0;  // 32'hc171311a;
    ram_cell[     459] = 32'h0;  // 32'he978ffe1;
    ram_cell[     460] = 32'h0;  // 32'h9cb806c0;
    ram_cell[     461] = 32'h0;  // 32'h9d20150e;
    ram_cell[     462] = 32'h0;  // 32'hf1df1e53;
    ram_cell[     463] = 32'h0;  // 32'h80cb3db7;
    ram_cell[     464] = 32'h0;  // 32'h71751e0b;
    ram_cell[     465] = 32'h0;  // 32'h01f0ed0c;
    ram_cell[     466] = 32'h0;  // 32'hba7fada6;
    ram_cell[     467] = 32'h0;  // 32'h966a6774;
    ram_cell[     468] = 32'h0;  // 32'h40857976;
    ram_cell[     469] = 32'h0;  // 32'h9b56987f;
    ram_cell[     470] = 32'h0;  // 32'hee4ad747;
    ram_cell[     471] = 32'h0;  // 32'h421fb8cd;
    ram_cell[     472] = 32'h0;  // 32'h47e1b407;
    ram_cell[     473] = 32'h0;  // 32'hd093c9e8;
    ram_cell[     474] = 32'h0;  // 32'hb6d05c0b;
    ram_cell[     475] = 32'h0;  // 32'h1f9017c2;
    ram_cell[     476] = 32'h0;  // 32'h3bebc027;
    ram_cell[     477] = 32'h0;  // 32'h804fa4f7;
    ram_cell[     478] = 32'h0;  // 32'ha5ed7407;
    ram_cell[     479] = 32'h0;  // 32'h92d57021;
    ram_cell[     480] = 32'h0;  // 32'h5440e8c4;
    ram_cell[     481] = 32'h0;  // 32'ha2d3bc68;
    ram_cell[     482] = 32'h0;  // 32'h6d2f3503;
    ram_cell[     483] = 32'h0;  // 32'h8f28d22b;
    ram_cell[     484] = 32'h0;  // 32'h88242010;
    ram_cell[     485] = 32'h0;  // 32'h7bebb632;
    ram_cell[     486] = 32'h0;  // 32'h0d8c3022;
    ram_cell[     487] = 32'h0;  // 32'h651754a1;
    ram_cell[     488] = 32'h0;  // 32'h676df589;
    ram_cell[     489] = 32'h0;  // 32'h6de6f6cd;
    ram_cell[     490] = 32'h0;  // 32'h62df79bc;
    ram_cell[     491] = 32'h0;  // 32'hea760de8;
    ram_cell[     492] = 32'h0;  // 32'hd4e11684;
    ram_cell[     493] = 32'h0;  // 32'h08d9bbd6;
    ram_cell[     494] = 32'h0;  // 32'haaa9fbc5;
    ram_cell[     495] = 32'h0;  // 32'h3bd3d918;
    ram_cell[     496] = 32'h0;  // 32'h1f9b4f78;
    ram_cell[     497] = 32'h0;  // 32'h8a026fbb;
    ram_cell[     498] = 32'h0;  // 32'h2fb929f6;
    ram_cell[     499] = 32'h0;  // 32'h83ccc770;
    ram_cell[     500] = 32'h0;  // 32'h974abe00;
    ram_cell[     501] = 32'h0;  // 32'h463e1b86;
    ram_cell[     502] = 32'h0;  // 32'h0413756f;
    ram_cell[     503] = 32'h0;  // 32'h17343dab;
    ram_cell[     504] = 32'h0;  // 32'h184b6e65;
    ram_cell[     505] = 32'h0;  // 32'he5e80ce1;
    ram_cell[     506] = 32'h0;  // 32'hdb218a5a;
    ram_cell[     507] = 32'h0;  // 32'haf4a0083;
    ram_cell[     508] = 32'h0;  // 32'h94c833fe;
    ram_cell[     509] = 32'h0;  // 32'hc163e695;
    ram_cell[     510] = 32'h0;  // 32'hccdf2993;
    ram_cell[     511] = 32'h0;  // 32'h74ea9752;
    ram_cell[     512] = 32'h0;  // 32'h5c49143f;
    ram_cell[     513] = 32'h0;  // 32'h4b0236e7;
    ram_cell[     514] = 32'h0;  // 32'hfecfbd41;
    ram_cell[     515] = 32'h0;  // 32'h0475c872;
    ram_cell[     516] = 32'h0;  // 32'h6d91be18;
    ram_cell[     517] = 32'h0;  // 32'hbea74503;
    ram_cell[     518] = 32'h0;  // 32'h2f4205da;
    ram_cell[     519] = 32'h0;  // 32'hc21c6c32;
    ram_cell[     520] = 32'h0;  // 32'hb6b462b1;
    ram_cell[     521] = 32'h0;  // 32'he7027dca;
    ram_cell[     522] = 32'h0;  // 32'h215b1553;
    ram_cell[     523] = 32'h0;  // 32'hbf2e22f8;
    ram_cell[     524] = 32'h0;  // 32'h73dc23f5;
    ram_cell[     525] = 32'h0;  // 32'hdc36f0a0;
    ram_cell[     526] = 32'h0;  // 32'h5fddedfd;
    ram_cell[     527] = 32'h0;  // 32'h00084891;
    ram_cell[     528] = 32'h0;  // 32'h1e03b36e;
    ram_cell[     529] = 32'h0;  // 32'h10dbcd82;
    ram_cell[     530] = 32'h0;  // 32'he63fe423;
    ram_cell[     531] = 32'h0;  // 32'h07964945;
    ram_cell[     532] = 32'h0;  // 32'h2d6e677f;
    ram_cell[     533] = 32'h0;  // 32'h852e8c60;
    ram_cell[     534] = 32'h0;  // 32'ha6a8babf;
    ram_cell[     535] = 32'h0;  // 32'h46a30fad;
    ram_cell[     536] = 32'h0;  // 32'h19d1b82c;
    ram_cell[     537] = 32'h0;  // 32'h98b70269;
    ram_cell[     538] = 32'h0;  // 32'hf88f74b1;
    ram_cell[     539] = 32'h0;  // 32'h95a64f00;
    ram_cell[     540] = 32'h0;  // 32'heb977522;
    ram_cell[     541] = 32'h0;  // 32'hae0775cc;
    ram_cell[     542] = 32'h0;  // 32'hf95699f9;
    ram_cell[     543] = 32'h0;  // 32'h1f2fc6c2;
    ram_cell[     544] = 32'h0;  // 32'hd44e524a;
    ram_cell[     545] = 32'h0;  // 32'h000ac059;
    ram_cell[     546] = 32'h0;  // 32'hed0439e8;
    ram_cell[     547] = 32'h0;  // 32'h22ad030e;
    ram_cell[     548] = 32'h0;  // 32'h902a423e;
    ram_cell[     549] = 32'h0;  // 32'h58059af3;
    ram_cell[     550] = 32'h0;  // 32'h855d9120;
    ram_cell[     551] = 32'h0;  // 32'h82ef96fb;
    ram_cell[     552] = 32'h0;  // 32'h33c8156a;
    ram_cell[     553] = 32'h0;  // 32'h4bc0a2cc;
    ram_cell[     554] = 32'h0;  // 32'heffb26e5;
    ram_cell[     555] = 32'h0;  // 32'h264e7821;
    ram_cell[     556] = 32'h0;  // 32'hb3145b89;
    ram_cell[     557] = 32'h0;  // 32'h9340a3b4;
    ram_cell[     558] = 32'h0;  // 32'h30e0e48f;
    ram_cell[     559] = 32'h0;  // 32'hafcdc14a;
    ram_cell[     560] = 32'h0;  // 32'haba9597f;
    ram_cell[     561] = 32'h0;  // 32'h55672fdd;
    ram_cell[     562] = 32'h0;  // 32'h708926f3;
    ram_cell[     563] = 32'h0;  // 32'h2b52eab5;
    ram_cell[     564] = 32'h0;  // 32'h40c646e3;
    ram_cell[     565] = 32'h0;  // 32'hf94ce171;
    ram_cell[     566] = 32'h0;  // 32'hdb6b4aa7;
    ram_cell[     567] = 32'h0;  // 32'h7f7b4d58;
    ram_cell[     568] = 32'h0;  // 32'h24b31f7d;
    ram_cell[     569] = 32'h0;  // 32'hc995bf22;
    ram_cell[     570] = 32'h0;  // 32'h21445fb0;
    ram_cell[     571] = 32'h0;  // 32'hce1655a3;
    ram_cell[     572] = 32'h0;  // 32'h7ba52c5f;
    ram_cell[     573] = 32'h0;  // 32'h88ceace9;
    ram_cell[     574] = 32'h0;  // 32'h37205130;
    ram_cell[     575] = 32'h0;  // 32'h3875bf48;
    ram_cell[     576] = 32'h0;  // 32'h09989464;
    ram_cell[     577] = 32'h0;  // 32'heb4a50cc;
    ram_cell[     578] = 32'h0;  // 32'h49d1081e;
    ram_cell[     579] = 32'h0;  // 32'hdb70831f;
    ram_cell[     580] = 32'h0;  // 32'hd3cf597c;
    ram_cell[     581] = 32'h0;  // 32'hf3096b38;
    ram_cell[     582] = 32'h0;  // 32'h260ac006;
    ram_cell[     583] = 32'h0;  // 32'h34b89c85;
    ram_cell[     584] = 32'h0;  // 32'h5dc0fa10;
    ram_cell[     585] = 32'h0;  // 32'h4814a6b1;
    ram_cell[     586] = 32'h0;  // 32'h43e5f795;
    ram_cell[     587] = 32'h0;  // 32'h9245ca3a;
    ram_cell[     588] = 32'h0;  // 32'hdc02c92c;
    ram_cell[     589] = 32'h0;  // 32'h2c7dcd16;
    ram_cell[     590] = 32'h0;  // 32'hf68239c7;
    ram_cell[     591] = 32'h0;  // 32'h3c3fc199;
    ram_cell[     592] = 32'h0;  // 32'h20ad6b8b;
    ram_cell[     593] = 32'h0;  // 32'hce307bc2;
    ram_cell[     594] = 32'h0;  // 32'h7ef3297d;
    ram_cell[     595] = 32'h0;  // 32'ha7cf2ef0;
    ram_cell[     596] = 32'h0;  // 32'h470be7ae;
    ram_cell[     597] = 32'h0;  // 32'h63e71d84;
    ram_cell[     598] = 32'h0;  // 32'h39d227b0;
    ram_cell[     599] = 32'h0;  // 32'h4119b8e7;
    ram_cell[     600] = 32'h0;  // 32'ha32cde97;
    ram_cell[     601] = 32'h0;  // 32'hd115832d;
    ram_cell[     602] = 32'h0;  // 32'hf9c9625c;
    ram_cell[     603] = 32'h0;  // 32'hd67dcc03;
    ram_cell[     604] = 32'h0;  // 32'h9b25c78d;
    ram_cell[     605] = 32'h0;  // 32'haef4aa84;
    ram_cell[     606] = 32'h0;  // 32'h8618d2f7;
    ram_cell[     607] = 32'h0;  // 32'h98547dbe;
    ram_cell[     608] = 32'h0;  // 32'hbf97c8f1;
    ram_cell[     609] = 32'h0;  // 32'h16ccef10;
    ram_cell[     610] = 32'h0;  // 32'hc78dda47;
    ram_cell[     611] = 32'h0;  // 32'h6bd6c19c;
    ram_cell[     612] = 32'h0;  // 32'hb3ffa756;
    ram_cell[     613] = 32'h0;  // 32'h13917058;
    ram_cell[     614] = 32'h0;  // 32'hd0078b89;
    ram_cell[     615] = 32'h0;  // 32'h3e2cdd6c;
    ram_cell[     616] = 32'h0;  // 32'h8ae4e8e1;
    ram_cell[     617] = 32'h0;  // 32'hada871b5;
    ram_cell[     618] = 32'h0;  // 32'hf6ee7c2a;
    ram_cell[     619] = 32'h0;  // 32'h41172310;
    ram_cell[     620] = 32'h0;  // 32'hf4ba1f15;
    ram_cell[     621] = 32'h0;  // 32'h7dac48da;
    ram_cell[     622] = 32'h0;  // 32'hd36961d0;
    ram_cell[     623] = 32'h0;  // 32'h2f90e55f;
    ram_cell[     624] = 32'h0;  // 32'h245638f3;
    ram_cell[     625] = 32'h0;  // 32'ha03d4dd2;
    ram_cell[     626] = 32'h0;  // 32'h8d8a99de;
    ram_cell[     627] = 32'h0;  // 32'h8608846b;
    ram_cell[     628] = 32'h0;  // 32'h1358bb09;
    ram_cell[     629] = 32'h0;  // 32'h2dc181d8;
    ram_cell[     630] = 32'h0;  // 32'h3cf093b8;
    ram_cell[     631] = 32'h0;  // 32'h94c1aa98;
    ram_cell[     632] = 32'h0;  // 32'h7896c028;
    ram_cell[     633] = 32'h0;  // 32'h18c4547d;
    ram_cell[     634] = 32'h0;  // 32'hd80d33ad;
    ram_cell[     635] = 32'h0;  // 32'h879baa13;
    ram_cell[     636] = 32'h0;  // 32'h0433e9e4;
    ram_cell[     637] = 32'h0;  // 32'h27e5019f;
    ram_cell[     638] = 32'h0;  // 32'hf5e4aded;
    ram_cell[     639] = 32'h0;  // 32'h9b3055f9;
    ram_cell[     640] = 32'h0;  // 32'h2ff74af7;
    ram_cell[     641] = 32'h0;  // 32'he950a18e;
    ram_cell[     642] = 32'h0;  // 32'h7d93f27a;
    ram_cell[     643] = 32'h0;  // 32'ha4905801;
    ram_cell[     644] = 32'h0;  // 32'ha3aaea8a;
    ram_cell[     645] = 32'h0;  // 32'h672f6dbf;
    ram_cell[     646] = 32'h0;  // 32'hf17aa7c8;
    ram_cell[     647] = 32'h0;  // 32'he14cfd85;
    ram_cell[     648] = 32'h0;  // 32'h6622b517;
    ram_cell[     649] = 32'h0;  // 32'h06d72c2a;
    ram_cell[     650] = 32'h0;  // 32'h7da36da0;
    ram_cell[     651] = 32'h0;  // 32'hdc6aee79;
    ram_cell[     652] = 32'h0;  // 32'h15cdf96f;
    ram_cell[     653] = 32'h0;  // 32'h075fab50;
    ram_cell[     654] = 32'h0;  // 32'h4884a45e;
    ram_cell[     655] = 32'h0;  // 32'hb97f6d26;
    ram_cell[     656] = 32'h0;  // 32'h19287063;
    ram_cell[     657] = 32'h0;  // 32'h576258d7;
    ram_cell[     658] = 32'h0;  // 32'h87e841ff;
    ram_cell[     659] = 32'h0;  // 32'ha856046f;
    ram_cell[     660] = 32'h0;  // 32'h2196bc26;
    ram_cell[     661] = 32'h0;  // 32'hbc059cab;
    ram_cell[     662] = 32'h0;  // 32'hdc712d53;
    ram_cell[     663] = 32'h0;  // 32'h7584d649;
    ram_cell[     664] = 32'h0;  // 32'h2238adf4;
    ram_cell[     665] = 32'h0;  // 32'hd9722f20;
    ram_cell[     666] = 32'h0;  // 32'h37c3e42f;
    ram_cell[     667] = 32'h0;  // 32'h6c832c25;
    ram_cell[     668] = 32'h0;  // 32'hdb3fc5a1;
    ram_cell[     669] = 32'h0;  // 32'h91d9924c;
    ram_cell[     670] = 32'h0;  // 32'hcf009b5a;
    ram_cell[     671] = 32'h0;  // 32'ha8ecdc56;
    ram_cell[     672] = 32'h0;  // 32'h5fb245b7;
    ram_cell[     673] = 32'h0;  // 32'hd02ed147;
    ram_cell[     674] = 32'h0;  // 32'h8fd3c5f2;
    ram_cell[     675] = 32'h0;  // 32'h99f6a6c2;
    ram_cell[     676] = 32'h0;  // 32'h8f17c8bf;
    ram_cell[     677] = 32'h0;  // 32'h46a5af3b;
    ram_cell[     678] = 32'h0;  // 32'hb0b1b32d;
    ram_cell[     679] = 32'h0;  // 32'h7ba82f53;
    ram_cell[     680] = 32'h0;  // 32'h89d821f5;
    ram_cell[     681] = 32'h0;  // 32'hca438b3f;
    ram_cell[     682] = 32'h0;  // 32'he50b7b97;
    ram_cell[     683] = 32'h0;  // 32'h759e8a3f;
    ram_cell[     684] = 32'h0;  // 32'h5e3dbf1b;
    ram_cell[     685] = 32'h0;  // 32'h8736675f;
    ram_cell[     686] = 32'h0;  // 32'hf76530de;
    ram_cell[     687] = 32'h0;  // 32'h4d85769d;
    ram_cell[     688] = 32'h0;  // 32'h2dbbe7a9;
    ram_cell[     689] = 32'h0;  // 32'h9d1ed4c4;
    ram_cell[     690] = 32'h0;  // 32'h8b99b936;
    ram_cell[     691] = 32'h0;  // 32'hb474157e;
    ram_cell[     692] = 32'h0;  // 32'hb52654dc;
    ram_cell[     693] = 32'h0;  // 32'h187ef830;
    ram_cell[     694] = 32'h0;  // 32'h60d9d566;
    ram_cell[     695] = 32'h0;  // 32'h2318eba6;
    ram_cell[     696] = 32'h0;  // 32'h575edec3;
    ram_cell[     697] = 32'h0;  // 32'hfe5adc7d;
    ram_cell[     698] = 32'h0;  // 32'ha5eead83;
    ram_cell[     699] = 32'h0;  // 32'h676e783e;
    ram_cell[     700] = 32'h0;  // 32'hccbfe1f2;
    ram_cell[     701] = 32'h0;  // 32'hc4d21366;
    ram_cell[     702] = 32'h0;  // 32'hfa0d4179;
    ram_cell[     703] = 32'h0;  // 32'h6081cf02;
    ram_cell[     704] = 32'h0;  // 32'h2fa17362;
    ram_cell[     705] = 32'h0;  // 32'h7a7952d2;
    ram_cell[     706] = 32'h0;  // 32'h88f199b3;
    ram_cell[     707] = 32'h0;  // 32'h6565fe84;
    ram_cell[     708] = 32'h0;  // 32'h382bceff;
    ram_cell[     709] = 32'h0;  // 32'h3d9c12d3;
    ram_cell[     710] = 32'h0;  // 32'h555a25b2;
    ram_cell[     711] = 32'h0;  // 32'h01a2af16;
    ram_cell[     712] = 32'h0;  // 32'h28a23b06;
    ram_cell[     713] = 32'h0;  // 32'hb484d067;
    ram_cell[     714] = 32'h0;  // 32'h37950be8;
    ram_cell[     715] = 32'h0;  // 32'h682233e4;
    ram_cell[     716] = 32'h0;  // 32'hf742f04e;
    ram_cell[     717] = 32'h0;  // 32'h8e0817a0;
    ram_cell[     718] = 32'h0;  // 32'hfe0ab0e5;
    ram_cell[     719] = 32'h0;  // 32'h1e3ca7af;
    ram_cell[     720] = 32'h0;  // 32'h5907540d;
    ram_cell[     721] = 32'h0;  // 32'hefe869a1;
    ram_cell[     722] = 32'h0;  // 32'h312962f7;
    ram_cell[     723] = 32'h0;  // 32'h1186f545;
    ram_cell[     724] = 32'h0;  // 32'h9be6004d;
    ram_cell[     725] = 32'h0;  // 32'h1b9674d7;
    ram_cell[     726] = 32'h0;  // 32'hfac35156;
    ram_cell[     727] = 32'h0;  // 32'ha238551f;
    ram_cell[     728] = 32'h0;  // 32'h662fb476;
    ram_cell[     729] = 32'h0;  // 32'hea773e4c;
    ram_cell[     730] = 32'h0;  // 32'h34f68238;
    ram_cell[     731] = 32'h0;  // 32'h19e60196;
    ram_cell[     732] = 32'h0;  // 32'h012dba64;
    ram_cell[     733] = 32'h0;  // 32'h439a2687;
    ram_cell[     734] = 32'h0;  // 32'hb5ad593b;
    ram_cell[     735] = 32'h0;  // 32'h11cae4f8;
    ram_cell[     736] = 32'h0;  // 32'h1079538f;
    ram_cell[     737] = 32'h0;  // 32'ha9fec724;
    ram_cell[     738] = 32'h0;  // 32'h4664b9b7;
    ram_cell[     739] = 32'h0;  // 32'hc8d102e7;
    ram_cell[     740] = 32'h0;  // 32'h85569387;
    ram_cell[     741] = 32'h0;  // 32'h32e4f282;
    ram_cell[     742] = 32'h0;  // 32'h15a8483f;
    ram_cell[     743] = 32'h0;  // 32'h8590d274;
    ram_cell[     744] = 32'h0;  // 32'h16f325ff;
    ram_cell[     745] = 32'h0;  // 32'h53ef4ac0;
    ram_cell[     746] = 32'h0;  // 32'hc63f325a;
    ram_cell[     747] = 32'h0;  // 32'h13e3012c;
    ram_cell[     748] = 32'h0;  // 32'h990ec75c;
    ram_cell[     749] = 32'h0;  // 32'h5c337435;
    ram_cell[     750] = 32'h0;  // 32'h0ad8cfb7;
    ram_cell[     751] = 32'h0;  // 32'h5914f8fa;
    ram_cell[     752] = 32'h0;  // 32'h1a53e98b;
    ram_cell[     753] = 32'h0;  // 32'hb6ccc8bc;
    ram_cell[     754] = 32'h0;  // 32'h25b197dd;
    ram_cell[     755] = 32'h0;  // 32'h0a86104c;
    ram_cell[     756] = 32'h0;  // 32'hd5e34854;
    ram_cell[     757] = 32'h0;  // 32'h77566d75;
    ram_cell[     758] = 32'h0;  // 32'h59330b82;
    ram_cell[     759] = 32'h0;  // 32'ha2e78e82;
    ram_cell[     760] = 32'h0;  // 32'h90b8d0e4;
    ram_cell[     761] = 32'h0;  // 32'he6f685d1;
    ram_cell[     762] = 32'h0;  // 32'h7d0a6727;
    ram_cell[     763] = 32'h0;  // 32'hc4839798;
    ram_cell[     764] = 32'h0;  // 32'h687742f5;
    ram_cell[     765] = 32'h0;  // 32'h60521638;
    ram_cell[     766] = 32'h0;  // 32'hef6cc205;
    ram_cell[     767] = 32'h0;  // 32'h82e76707;
    ram_cell[     768] = 32'h0;  // 32'h20d09c6a;
    ram_cell[     769] = 32'h0;  // 32'h5c4cd756;
    ram_cell[     770] = 32'h0;  // 32'ha26d6852;
    ram_cell[     771] = 32'h0;  // 32'h1aa9ea73;
    ram_cell[     772] = 32'h0;  // 32'h9ebe227c;
    ram_cell[     773] = 32'h0;  // 32'hbecf27ed;
    ram_cell[     774] = 32'h0;  // 32'hb73d231f;
    ram_cell[     775] = 32'h0;  // 32'hd9826d13;
    ram_cell[     776] = 32'h0;  // 32'hf2dd9dee;
    ram_cell[     777] = 32'h0;  // 32'h324c2a15;
    ram_cell[     778] = 32'h0;  // 32'hc9ad294e;
    ram_cell[     779] = 32'h0;  // 32'hc07c878f;
    ram_cell[     780] = 32'h0;  // 32'h47ff1742;
    ram_cell[     781] = 32'h0;  // 32'hf78dd6ae;
    ram_cell[     782] = 32'h0;  // 32'h436489d9;
    ram_cell[     783] = 32'h0;  // 32'h80ca423c;
    ram_cell[     784] = 32'h0;  // 32'hc24dcaaf;
    ram_cell[     785] = 32'h0;  // 32'h9d9650c3;
    ram_cell[     786] = 32'h0;  // 32'h7b59baeb;
    ram_cell[     787] = 32'h0;  // 32'h593f8a01;
    ram_cell[     788] = 32'h0;  // 32'h0a5de71b;
    ram_cell[     789] = 32'h0;  // 32'hbacda91c;
    ram_cell[     790] = 32'h0;  // 32'h11449961;
    ram_cell[     791] = 32'h0;  // 32'h8556fbb1;
    ram_cell[     792] = 32'h0;  // 32'h808abc4e;
    ram_cell[     793] = 32'h0;  // 32'h98530c31;
    ram_cell[     794] = 32'h0;  // 32'hed8530fc;
    ram_cell[     795] = 32'h0;  // 32'h6c3d7698;
    ram_cell[     796] = 32'h0;  // 32'hd8ebd6ef;
    ram_cell[     797] = 32'h0;  // 32'hb9d6174c;
    ram_cell[     798] = 32'h0;  // 32'h7d466ab9;
    ram_cell[     799] = 32'h0;  // 32'hc2f70e4a;
    ram_cell[     800] = 32'h0;  // 32'h9d6d9ca6;
    ram_cell[     801] = 32'h0;  // 32'ha29a7d2a;
    ram_cell[     802] = 32'h0;  // 32'heb67095a;
    ram_cell[     803] = 32'h0;  // 32'h01033857;
    ram_cell[     804] = 32'h0;  // 32'ha66a190c;
    ram_cell[     805] = 32'h0;  // 32'he7e9aa9a;
    ram_cell[     806] = 32'h0;  // 32'h1bc284d6;
    ram_cell[     807] = 32'h0;  // 32'hc71ef6e6;
    ram_cell[     808] = 32'h0;  // 32'ha11581a8;
    ram_cell[     809] = 32'h0;  // 32'hb4f93b7f;
    ram_cell[     810] = 32'h0;  // 32'hef6762e0;
    ram_cell[     811] = 32'h0;  // 32'h26616ec8;
    ram_cell[     812] = 32'h0;  // 32'h47287838;
    ram_cell[     813] = 32'h0;  // 32'h252d4dd6;
    ram_cell[     814] = 32'h0;  // 32'h051fc8b3;
    ram_cell[     815] = 32'h0;  // 32'hd1cf16ea;
    ram_cell[     816] = 32'h0;  // 32'h57ccc258;
    ram_cell[     817] = 32'h0;  // 32'h4007d8d9;
    ram_cell[     818] = 32'h0;  // 32'hd3e945e7;
    ram_cell[     819] = 32'h0;  // 32'h542eb391;
    ram_cell[     820] = 32'h0;  // 32'h899411d5;
    ram_cell[     821] = 32'h0;  // 32'haca5ae17;
    ram_cell[     822] = 32'h0;  // 32'h2fb99992;
    ram_cell[     823] = 32'h0;  // 32'hff0d2248;
    ram_cell[     824] = 32'h0;  // 32'h71e983ce;
    ram_cell[     825] = 32'h0;  // 32'he8e49bfc;
    ram_cell[     826] = 32'h0;  // 32'h8443263a;
    ram_cell[     827] = 32'h0;  // 32'h91072ca4;
    ram_cell[     828] = 32'h0;  // 32'hc5d9e07e;
    ram_cell[     829] = 32'h0;  // 32'hcf90efeb;
    ram_cell[     830] = 32'h0;  // 32'ha6e12f10;
    ram_cell[     831] = 32'h0;  // 32'he7897735;
    ram_cell[     832] = 32'h0;  // 32'h1f83704b;
    ram_cell[     833] = 32'h0;  // 32'hcd637447;
    ram_cell[     834] = 32'h0;  // 32'h68c8f71c;
    ram_cell[     835] = 32'h0;  // 32'hd1e3289a;
    ram_cell[     836] = 32'h0;  // 32'hd80957c4;
    ram_cell[     837] = 32'h0;  // 32'hf17d900c;
    ram_cell[     838] = 32'h0;  // 32'h18347f58;
    ram_cell[     839] = 32'h0;  // 32'hedfb93d8;
    ram_cell[     840] = 32'h0;  // 32'h01c1cda9;
    ram_cell[     841] = 32'h0;  // 32'hb56a8bef;
    ram_cell[     842] = 32'h0;  // 32'hca0de49a;
    ram_cell[     843] = 32'h0;  // 32'hf0710b14;
    ram_cell[     844] = 32'h0;  // 32'h573c75b1;
    ram_cell[     845] = 32'h0;  // 32'h058c0a78;
    ram_cell[     846] = 32'h0;  // 32'h11398b86;
    ram_cell[     847] = 32'h0;  // 32'ha6d12d03;
    ram_cell[     848] = 32'h0;  // 32'hafc85fe2;
    ram_cell[     849] = 32'h0;  // 32'h82f51fc5;
    ram_cell[     850] = 32'h0;  // 32'hc7ce7230;
    ram_cell[     851] = 32'h0;  // 32'h10524f79;
    ram_cell[     852] = 32'h0;  // 32'hb70f8665;
    ram_cell[     853] = 32'h0;  // 32'h2125d40e;
    ram_cell[     854] = 32'h0;  // 32'h21c6a074;
    ram_cell[     855] = 32'h0;  // 32'h19c13ae1;
    ram_cell[     856] = 32'h0;  // 32'h846c2436;
    ram_cell[     857] = 32'h0;  // 32'h27334b11;
    ram_cell[     858] = 32'h0;  // 32'h1994b115;
    ram_cell[     859] = 32'h0;  // 32'h26f37d5b;
    ram_cell[     860] = 32'h0;  // 32'h78b2a1d1;
    ram_cell[     861] = 32'h0;  // 32'h9e831e0f;
    ram_cell[     862] = 32'h0;  // 32'hb95b5161;
    ram_cell[     863] = 32'h0;  // 32'hfc431c2e;
    ram_cell[     864] = 32'h0;  // 32'h7e5cd301;
    ram_cell[     865] = 32'h0;  // 32'h4e2f2d30;
    ram_cell[     866] = 32'h0;  // 32'haacdd442;
    ram_cell[     867] = 32'h0;  // 32'h564aefc6;
    ram_cell[     868] = 32'h0;  // 32'hd966c107;
    ram_cell[     869] = 32'h0;  // 32'h4e502a06;
    ram_cell[     870] = 32'h0;  // 32'h833424a3;
    ram_cell[     871] = 32'h0;  // 32'hcc678c56;
    ram_cell[     872] = 32'h0;  // 32'hc752a951;
    ram_cell[     873] = 32'h0;  // 32'hd73ed4fc;
    ram_cell[     874] = 32'h0;  // 32'hee1e967a;
    ram_cell[     875] = 32'h0;  // 32'h6b307543;
    ram_cell[     876] = 32'h0;  // 32'h021d7c8c;
    ram_cell[     877] = 32'h0;  // 32'ha88b49ea;
    ram_cell[     878] = 32'h0;  // 32'h51d03186;
    ram_cell[     879] = 32'h0;  // 32'h2e508f1a;
    ram_cell[     880] = 32'h0;  // 32'h01671dfc;
    ram_cell[     881] = 32'h0;  // 32'hd1e9a60e;
    ram_cell[     882] = 32'h0;  // 32'hf32e2448;
    ram_cell[     883] = 32'h0;  // 32'h9ca094e9;
    ram_cell[     884] = 32'h0;  // 32'h8ad7e460;
    ram_cell[     885] = 32'h0;  // 32'h3eaea1d5;
    ram_cell[     886] = 32'h0;  // 32'h9e891184;
    ram_cell[     887] = 32'h0;  // 32'h2fe32e25;
    ram_cell[     888] = 32'h0;  // 32'hce74e9fb;
    ram_cell[     889] = 32'h0;  // 32'h6708179c;
    ram_cell[     890] = 32'h0;  // 32'h8128ba2b;
    ram_cell[     891] = 32'h0;  // 32'h5c16b2b1;
    ram_cell[     892] = 32'h0;  // 32'h18b087b4;
    ram_cell[     893] = 32'h0;  // 32'had1dddf5;
    ram_cell[     894] = 32'h0;  // 32'h70bae58e;
    ram_cell[     895] = 32'h0;  // 32'h5979c6ee;
    ram_cell[     896] = 32'h0;  // 32'h94ab2060;
    ram_cell[     897] = 32'h0;  // 32'h2726bc53;
    ram_cell[     898] = 32'h0;  // 32'h8c1c253e;
    ram_cell[     899] = 32'h0;  // 32'h14c5f81d;
    ram_cell[     900] = 32'h0;  // 32'ha9e846c0;
    ram_cell[     901] = 32'h0;  // 32'h2529fc99;
    ram_cell[     902] = 32'h0;  // 32'hdc5ee4cf;
    ram_cell[     903] = 32'h0;  // 32'hed65a638;
    ram_cell[     904] = 32'h0;  // 32'ha58df84e;
    ram_cell[     905] = 32'h0;  // 32'h3d7b5c2c;
    ram_cell[     906] = 32'h0;  // 32'hee1bb5f8;
    ram_cell[     907] = 32'h0;  // 32'hae131489;
    ram_cell[     908] = 32'h0;  // 32'h13549384;
    ram_cell[     909] = 32'h0;  // 32'h49bea1c7;
    ram_cell[     910] = 32'h0;  // 32'h9d5f8761;
    ram_cell[     911] = 32'h0;  // 32'h1d3fa6c2;
    ram_cell[     912] = 32'h0;  // 32'h54800a8e;
    ram_cell[     913] = 32'h0;  // 32'h1f6a960d;
    ram_cell[     914] = 32'h0;  // 32'h8e8c82cb;
    ram_cell[     915] = 32'h0;  // 32'h9f641846;
    ram_cell[     916] = 32'h0;  // 32'hedacd512;
    ram_cell[     917] = 32'h0;  // 32'h212dbe42;
    ram_cell[     918] = 32'h0;  // 32'h14c33429;
    ram_cell[     919] = 32'h0;  // 32'hdf5507ca;
    ram_cell[     920] = 32'h0;  // 32'h9649ce90;
    ram_cell[     921] = 32'h0;  // 32'h8455e365;
    ram_cell[     922] = 32'h0;  // 32'h64574965;
    ram_cell[     923] = 32'h0;  // 32'h45f4746b;
    ram_cell[     924] = 32'h0;  // 32'h211a2851;
    ram_cell[     925] = 32'h0;  // 32'h081ba044;
    ram_cell[     926] = 32'h0;  // 32'hc717ac58;
    ram_cell[     927] = 32'h0;  // 32'h4a6e49ca;
    ram_cell[     928] = 32'h0;  // 32'h4b2c86b5;
    ram_cell[     929] = 32'h0;  // 32'h688f7a68;
    ram_cell[     930] = 32'h0;  // 32'h58bad1fe;
    ram_cell[     931] = 32'h0;  // 32'h0a0341be;
    ram_cell[     932] = 32'h0;  // 32'h80fbff7d;
    ram_cell[     933] = 32'h0;  // 32'hdba5ab07;
    ram_cell[     934] = 32'h0;  // 32'h0f6ceeb0;
    ram_cell[     935] = 32'h0;  // 32'he3c53a10;
    ram_cell[     936] = 32'h0;  // 32'hd24e5eb4;
    ram_cell[     937] = 32'h0;  // 32'h5726e76d;
    ram_cell[     938] = 32'h0;  // 32'hc803d836;
    ram_cell[     939] = 32'h0;  // 32'he47d250b;
    ram_cell[     940] = 32'h0;  // 32'hc522edf4;
    ram_cell[     941] = 32'h0;  // 32'h07baad6f;
    ram_cell[     942] = 32'h0;  // 32'hbc35d114;
    ram_cell[     943] = 32'h0;  // 32'h1ce1f0ea;
    ram_cell[     944] = 32'h0;  // 32'h49d9adfe;
    ram_cell[     945] = 32'h0;  // 32'he5bfd913;
    ram_cell[     946] = 32'h0;  // 32'h0b74f4d3;
    ram_cell[     947] = 32'h0;  // 32'h27a53d5a;
    ram_cell[     948] = 32'h0;  // 32'h1e251c98;
    ram_cell[     949] = 32'h0;  // 32'h9f803a39;
    ram_cell[     950] = 32'h0;  // 32'h33b3c529;
    ram_cell[     951] = 32'h0;  // 32'ha2010851;
    ram_cell[     952] = 32'h0;  // 32'h7b207b30;
    ram_cell[     953] = 32'h0;  // 32'h8854d44a;
    ram_cell[     954] = 32'h0;  // 32'h2de59c89;
    ram_cell[     955] = 32'h0;  // 32'hb51c6a23;
    ram_cell[     956] = 32'h0;  // 32'hf9f3a81e;
    ram_cell[     957] = 32'h0;  // 32'h5f2c048f;
    ram_cell[     958] = 32'h0;  // 32'hf1d2886b;
    ram_cell[     959] = 32'h0;  // 32'h6fc187e1;
    ram_cell[     960] = 32'h0;  // 32'h8343ad28;
    ram_cell[     961] = 32'h0;  // 32'h941eeb94;
    ram_cell[     962] = 32'h0;  // 32'h88fe668c;
    ram_cell[     963] = 32'h0;  // 32'hd9e0756a;
    ram_cell[     964] = 32'h0;  // 32'h2b61bb21;
    ram_cell[     965] = 32'h0;  // 32'he60fe1b8;
    ram_cell[     966] = 32'h0;  // 32'h03848404;
    ram_cell[     967] = 32'h0;  // 32'h6007589e;
    ram_cell[     968] = 32'h0;  // 32'h9ef8846c;
    ram_cell[     969] = 32'h0;  // 32'h3cbca4da;
    ram_cell[     970] = 32'h0;  // 32'he325306f;
    ram_cell[     971] = 32'h0;  // 32'hca1aa03d;
    ram_cell[     972] = 32'h0;  // 32'h4b0d628c;
    ram_cell[     973] = 32'h0;  // 32'h31f5ac0c;
    ram_cell[     974] = 32'h0;  // 32'h86cf93a5;
    ram_cell[     975] = 32'h0;  // 32'hac24c8cb;
    ram_cell[     976] = 32'h0;  // 32'he502f603;
    ram_cell[     977] = 32'h0;  // 32'hf8886804;
    ram_cell[     978] = 32'h0;  // 32'hca39feae;
    ram_cell[     979] = 32'h0;  // 32'h4b1fd1e3;
    ram_cell[     980] = 32'h0;  // 32'h21739904;
    ram_cell[     981] = 32'h0;  // 32'he16fad27;
    ram_cell[     982] = 32'h0;  // 32'hd4d04917;
    ram_cell[     983] = 32'h0;  // 32'h47fb521d;
    ram_cell[     984] = 32'h0;  // 32'hf3b25edc;
    ram_cell[     985] = 32'h0;  // 32'h8ed2a284;
    ram_cell[     986] = 32'h0;  // 32'hc0eb20d4;
    ram_cell[     987] = 32'h0;  // 32'h87110f82;
    ram_cell[     988] = 32'h0;  // 32'h68e4bf1a;
    ram_cell[     989] = 32'h0;  // 32'hb9d9e51a;
    ram_cell[     990] = 32'h0;  // 32'hb7cd69c4;
    ram_cell[     991] = 32'h0;  // 32'h37f5417b;
    ram_cell[     992] = 32'h0;  // 32'hfb33754d;
    ram_cell[     993] = 32'h0;  // 32'h36c6f78c;
    ram_cell[     994] = 32'h0;  // 32'hca7c55fb;
    ram_cell[     995] = 32'h0;  // 32'h7cdefb49;
    ram_cell[     996] = 32'h0;  // 32'h23d4b2e6;
    ram_cell[     997] = 32'h0;  // 32'hc05af670;
    ram_cell[     998] = 32'h0;  // 32'h4192b675;
    ram_cell[     999] = 32'h0;  // 32'h232e55d0;
    ram_cell[    1000] = 32'h0;  // 32'h8f133c61;
    ram_cell[    1001] = 32'h0;  // 32'h2770a16a;
    ram_cell[    1002] = 32'h0;  // 32'hf7df8b11;
    ram_cell[    1003] = 32'h0;  // 32'hb9dab935;
    ram_cell[    1004] = 32'h0;  // 32'h051a1053;
    ram_cell[    1005] = 32'h0;  // 32'h9dbc0518;
    ram_cell[    1006] = 32'h0;  // 32'h81a95dbb;
    ram_cell[    1007] = 32'h0;  // 32'hac59e164;
    ram_cell[    1008] = 32'h0;  // 32'h9cfde310;
    ram_cell[    1009] = 32'h0;  // 32'h1cc152f7;
    ram_cell[    1010] = 32'h0;  // 32'h2c0fe90d;
    ram_cell[    1011] = 32'h0;  // 32'hc9a3536b;
    ram_cell[    1012] = 32'h0;  // 32'h74cb7558;
    ram_cell[    1013] = 32'h0;  // 32'h812d328f;
    ram_cell[    1014] = 32'h0;  // 32'h088dd765;
    ram_cell[    1015] = 32'h0;  // 32'h188aabbd;
    ram_cell[    1016] = 32'h0;  // 32'hfe85b606;
    ram_cell[    1017] = 32'h0;  // 32'h61dbd168;
    ram_cell[    1018] = 32'h0;  // 32'h89c7f1af;
    ram_cell[    1019] = 32'h0;  // 32'hb2846959;
    ram_cell[    1020] = 32'h0;  // 32'h000dbf76;
    ram_cell[    1021] = 32'h0;  // 32'ha280d3dd;
    ram_cell[    1022] = 32'h0;  // 32'h5615b9de;
    ram_cell[    1023] = 32'h0;  // 32'hf09eefd2;
    // src matrix A
    ram_cell[    1024] = 32'h3ac28bc9;
    ram_cell[    1025] = 32'h21d990cf;
    ram_cell[    1026] = 32'h2477ae53;
    ram_cell[    1027] = 32'hddff7972;
    ram_cell[    1028] = 32'hbfc842ed;
    ram_cell[    1029] = 32'hae9718cb;
    ram_cell[    1030] = 32'hf96e3497;
    ram_cell[    1031] = 32'hd165382f;
    ram_cell[    1032] = 32'h3c948d30;
    ram_cell[    1033] = 32'h137f41c4;
    ram_cell[    1034] = 32'h085809ad;
    ram_cell[    1035] = 32'h4f072c1d;
    ram_cell[    1036] = 32'hb3664c63;
    ram_cell[    1037] = 32'h295ee0d6;
    ram_cell[    1038] = 32'hf70d4879;
    ram_cell[    1039] = 32'h9c61747e;
    ram_cell[    1040] = 32'h965c5a61;
    ram_cell[    1041] = 32'h8a8e09d0;
    ram_cell[    1042] = 32'h4e401610;
    ram_cell[    1043] = 32'hc4348f08;
    ram_cell[    1044] = 32'hbaba2803;
    ram_cell[    1045] = 32'h489cea69;
    ram_cell[    1046] = 32'h19854cd6;
    ram_cell[    1047] = 32'h657eb168;
    ram_cell[    1048] = 32'h7b9f5af2;
    ram_cell[    1049] = 32'h9dab7c28;
    ram_cell[    1050] = 32'hcb32bc6b;
    ram_cell[    1051] = 32'hf9f676ef;
    ram_cell[    1052] = 32'h2ac78c29;
    ram_cell[    1053] = 32'hdee1d521;
    ram_cell[    1054] = 32'h188fd936;
    ram_cell[    1055] = 32'ha50197aa;
    ram_cell[    1056] = 32'h09b1bf9e;
    ram_cell[    1057] = 32'h7f808656;
    ram_cell[    1058] = 32'he3a48c30;
    ram_cell[    1059] = 32'haefcc162;
    ram_cell[    1060] = 32'h72939a4b;
    ram_cell[    1061] = 32'h972d0f18;
    ram_cell[    1062] = 32'hada11242;
    ram_cell[    1063] = 32'he4e89550;
    ram_cell[    1064] = 32'h4e377177;
    ram_cell[    1065] = 32'hf9ab0e2b;
    ram_cell[    1066] = 32'hb2204add;
    ram_cell[    1067] = 32'h3f495ac6;
    ram_cell[    1068] = 32'h7bd83270;
    ram_cell[    1069] = 32'h0db82cd2;
    ram_cell[    1070] = 32'hf321b534;
    ram_cell[    1071] = 32'had3a17bc;
    ram_cell[    1072] = 32'hfce4c176;
    ram_cell[    1073] = 32'hf245620a;
    ram_cell[    1074] = 32'h403734cb;
    ram_cell[    1075] = 32'h12523322;
    ram_cell[    1076] = 32'h232c4ddd;
    ram_cell[    1077] = 32'h40690188;
    ram_cell[    1078] = 32'haa3cc187;
    ram_cell[    1079] = 32'h07468e21;
    ram_cell[    1080] = 32'hf56eac69;
    ram_cell[    1081] = 32'ha9e8e7f5;
    ram_cell[    1082] = 32'h5802c8fb;
    ram_cell[    1083] = 32'hac35edc0;
    ram_cell[    1084] = 32'hceb1dfdb;
    ram_cell[    1085] = 32'h31d441fc;
    ram_cell[    1086] = 32'h3360df0c;
    ram_cell[    1087] = 32'h6d8557b5;
    ram_cell[    1088] = 32'hfffcdafd;
    ram_cell[    1089] = 32'h30c3cd9f;
    ram_cell[    1090] = 32'hee876d20;
    ram_cell[    1091] = 32'h795be524;
    ram_cell[    1092] = 32'h23f33cf4;
    ram_cell[    1093] = 32'h022cc3fc;
    ram_cell[    1094] = 32'h0baa7f7b;
    ram_cell[    1095] = 32'h81b72ad2;
    ram_cell[    1096] = 32'h470e33a3;
    ram_cell[    1097] = 32'h506c6730;
    ram_cell[    1098] = 32'h8e8ba40b;
    ram_cell[    1099] = 32'h93f4feea;
    ram_cell[    1100] = 32'hbde56566;
    ram_cell[    1101] = 32'h867e3960;
    ram_cell[    1102] = 32'ha7f596bb;
    ram_cell[    1103] = 32'hc02100f0;
    ram_cell[    1104] = 32'hcdb46e17;
    ram_cell[    1105] = 32'hf01dd821;
    ram_cell[    1106] = 32'h0506d6d7;
    ram_cell[    1107] = 32'hacd165fa;
    ram_cell[    1108] = 32'h8b8be1e5;
    ram_cell[    1109] = 32'hba154db6;
    ram_cell[    1110] = 32'h510be11b;
    ram_cell[    1111] = 32'hbe207165;
    ram_cell[    1112] = 32'hd50aaeab;
    ram_cell[    1113] = 32'h95a30f29;
    ram_cell[    1114] = 32'ha3d17ccf;
    ram_cell[    1115] = 32'h4452bdf5;
    ram_cell[    1116] = 32'hfaee4d95;
    ram_cell[    1117] = 32'hce1b7bbb;
    ram_cell[    1118] = 32'h31fa5e2c;
    ram_cell[    1119] = 32'h4c83b65f;
    ram_cell[    1120] = 32'h6097d60c;
    ram_cell[    1121] = 32'h7de19fa7;
    ram_cell[    1122] = 32'h0187ac9d;
    ram_cell[    1123] = 32'h7557fb7d;
    ram_cell[    1124] = 32'h395dff9b;
    ram_cell[    1125] = 32'hd978d73b;
    ram_cell[    1126] = 32'h0da20b20;
    ram_cell[    1127] = 32'hccdd0953;
    ram_cell[    1128] = 32'ha84180a6;
    ram_cell[    1129] = 32'hc000041b;
    ram_cell[    1130] = 32'hf5867791;
    ram_cell[    1131] = 32'h6f8ff3e1;
    ram_cell[    1132] = 32'h9828ed73;
    ram_cell[    1133] = 32'hd0f3d12f;
    ram_cell[    1134] = 32'h62e2d177;
    ram_cell[    1135] = 32'h2260fd9b;
    ram_cell[    1136] = 32'h0bf1768b;
    ram_cell[    1137] = 32'h390ee726;
    ram_cell[    1138] = 32'hefb4c525;
    ram_cell[    1139] = 32'h8de61b34;
    ram_cell[    1140] = 32'h81788219;
    ram_cell[    1141] = 32'he75069b0;
    ram_cell[    1142] = 32'hfbe5cbe7;
    ram_cell[    1143] = 32'he9d2f0ca;
    ram_cell[    1144] = 32'h9b631958;
    ram_cell[    1145] = 32'h18be72fd;
    ram_cell[    1146] = 32'h483501c2;
    ram_cell[    1147] = 32'h57a3f038;
    ram_cell[    1148] = 32'he0f4e809;
    ram_cell[    1149] = 32'h62344722;
    ram_cell[    1150] = 32'h2d660e0c;
    ram_cell[    1151] = 32'h1e4ba66a;
    ram_cell[    1152] = 32'h85d84aa1;
    ram_cell[    1153] = 32'h918bd820;
    ram_cell[    1154] = 32'hbbd3f1d4;
    ram_cell[    1155] = 32'h75fbad06;
    ram_cell[    1156] = 32'h4ee43c8e;
    ram_cell[    1157] = 32'h54480eac;
    ram_cell[    1158] = 32'h3b041e70;
    ram_cell[    1159] = 32'h1a4f77ce;
    ram_cell[    1160] = 32'h58b388a8;
    ram_cell[    1161] = 32'had3628c4;
    ram_cell[    1162] = 32'h9fb0e0fc;
    ram_cell[    1163] = 32'h92ffb3bc;
    ram_cell[    1164] = 32'hec1360a0;
    ram_cell[    1165] = 32'hd2ce3d1f;
    ram_cell[    1166] = 32'h1cc71801;
    ram_cell[    1167] = 32'h23246d0f;
    ram_cell[    1168] = 32'h5ee713d3;
    ram_cell[    1169] = 32'h11462ffb;
    ram_cell[    1170] = 32'h59724695;
    ram_cell[    1171] = 32'h0c3588e4;
    ram_cell[    1172] = 32'h473b5d0b;
    ram_cell[    1173] = 32'hba5a18e1;
    ram_cell[    1174] = 32'h94992f57;
    ram_cell[    1175] = 32'ha602b74e;
    ram_cell[    1176] = 32'h5ca4228f;
    ram_cell[    1177] = 32'h793bddc1;
    ram_cell[    1178] = 32'h2758f665;
    ram_cell[    1179] = 32'h5f8ed1e4;
    ram_cell[    1180] = 32'h8db9a6f0;
    ram_cell[    1181] = 32'h25557194;
    ram_cell[    1182] = 32'h9718a6a2;
    ram_cell[    1183] = 32'h1e1df912;
    ram_cell[    1184] = 32'ha9b3eb3a;
    ram_cell[    1185] = 32'h7ff83303;
    ram_cell[    1186] = 32'h91691dd1;
    ram_cell[    1187] = 32'h4731254a;
    ram_cell[    1188] = 32'ha8ae9540;
    ram_cell[    1189] = 32'h3d78c1c8;
    ram_cell[    1190] = 32'h6c1c4eeb;
    ram_cell[    1191] = 32'he59c301c;
    ram_cell[    1192] = 32'hbedc9f0d;
    ram_cell[    1193] = 32'h3ce4cda8;
    ram_cell[    1194] = 32'h0a6e3e44;
    ram_cell[    1195] = 32'h8ad20403;
    ram_cell[    1196] = 32'h116220f0;
    ram_cell[    1197] = 32'h662c3513;
    ram_cell[    1198] = 32'h1b6951a7;
    ram_cell[    1199] = 32'h4d04fe7a;
    ram_cell[    1200] = 32'hdd0bfe87;
    ram_cell[    1201] = 32'h4710a8a5;
    ram_cell[    1202] = 32'h34fc53f4;
    ram_cell[    1203] = 32'h9ad03dd2;
    ram_cell[    1204] = 32'hfd59a538;
    ram_cell[    1205] = 32'h5d578a18;
    ram_cell[    1206] = 32'h6fae8dcb;
    ram_cell[    1207] = 32'h2a73d021;
    ram_cell[    1208] = 32'h7b6935df;
    ram_cell[    1209] = 32'h25298f64;
    ram_cell[    1210] = 32'h2a900edb;
    ram_cell[    1211] = 32'h2655892f;
    ram_cell[    1212] = 32'h83ded03a;
    ram_cell[    1213] = 32'h84524b4e;
    ram_cell[    1214] = 32'he3873e77;
    ram_cell[    1215] = 32'hea70043b;
    ram_cell[    1216] = 32'ha5d3ec5d;
    ram_cell[    1217] = 32'h4893ccc7;
    ram_cell[    1218] = 32'hbdf93b77;
    ram_cell[    1219] = 32'h39ccc5d6;
    ram_cell[    1220] = 32'h7291d459;
    ram_cell[    1221] = 32'h99996564;
    ram_cell[    1222] = 32'hde98f990;
    ram_cell[    1223] = 32'h3cb008e8;
    ram_cell[    1224] = 32'h4e074994;
    ram_cell[    1225] = 32'hf573a78f;
    ram_cell[    1226] = 32'h0511ebaf;
    ram_cell[    1227] = 32'h85dabf5b;
    ram_cell[    1228] = 32'h5e7089a0;
    ram_cell[    1229] = 32'h45e2b7c8;
    ram_cell[    1230] = 32'h30781c3d;
    ram_cell[    1231] = 32'hb144cf59;
    ram_cell[    1232] = 32'h8e20cc8a;
    ram_cell[    1233] = 32'h5bc8a72a;
    ram_cell[    1234] = 32'hd491bef4;
    ram_cell[    1235] = 32'h5d342a90;
    ram_cell[    1236] = 32'h961d27d3;
    ram_cell[    1237] = 32'h1348914c;
    ram_cell[    1238] = 32'h663fe6b0;
    ram_cell[    1239] = 32'he75afd52;
    ram_cell[    1240] = 32'h3b5ebf58;
    ram_cell[    1241] = 32'he363c1fb;
    ram_cell[    1242] = 32'h7c2caf1f;
    ram_cell[    1243] = 32'h58f7b35a;
    ram_cell[    1244] = 32'h340b26e0;
    ram_cell[    1245] = 32'h31b24bba;
    ram_cell[    1246] = 32'h80bf8214;
    ram_cell[    1247] = 32'h8ba382d8;
    ram_cell[    1248] = 32'h0d81fd4c;
    ram_cell[    1249] = 32'h4547925d;
    ram_cell[    1250] = 32'h545eac18;
    ram_cell[    1251] = 32'hf9424417;
    ram_cell[    1252] = 32'he3aaac6a;
    ram_cell[    1253] = 32'h0fefa1a0;
    ram_cell[    1254] = 32'hc0fe760a;
    ram_cell[    1255] = 32'hf291bfe0;
    ram_cell[    1256] = 32'h27fca090;
    ram_cell[    1257] = 32'he3689743;
    ram_cell[    1258] = 32'h6fd33f56;
    ram_cell[    1259] = 32'h1517a5dc;
    ram_cell[    1260] = 32'hef932823;
    ram_cell[    1261] = 32'heda6df5a;
    ram_cell[    1262] = 32'heee14924;
    ram_cell[    1263] = 32'h49d851f6;
    ram_cell[    1264] = 32'h433f3ae0;
    ram_cell[    1265] = 32'h7742fd9b;
    ram_cell[    1266] = 32'h5fdf00ea;
    ram_cell[    1267] = 32'h2a508e64;
    ram_cell[    1268] = 32'h3f8714d3;
    ram_cell[    1269] = 32'h78c43fa4;
    ram_cell[    1270] = 32'hd9f22ac8;
    ram_cell[    1271] = 32'h919195fe;
    ram_cell[    1272] = 32'h4bce79d7;
    ram_cell[    1273] = 32'ha0b370c8;
    ram_cell[    1274] = 32'h17ecabbf;
    ram_cell[    1275] = 32'h6f76a232;
    ram_cell[    1276] = 32'hd60abec8;
    ram_cell[    1277] = 32'h7133f073;
    ram_cell[    1278] = 32'h9ef94d53;
    ram_cell[    1279] = 32'h69ae12a3;
    ram_cell[    1280] = 32'ha51d556b;
    ram_cell[    1281] = 32'h6f90670d;
    ram_cell[    1282] = 32'hf6f5eaa8;
    ram_cell[    1283] = 32'hffc63da6;
    ram_cell[    1284] = 32'h6bf4ac52;
    ram_cell[    1285] = 32'hb0083aa3;
    ram_cell[    1286] = 32'h6046ab89;
    ram_cell[    1287] = 32'h11929dc2;
    ram_cell[    1288] = 32'hc08311d8;
    ram_cell[    1289] = 32'h87c13d6a;
    ram_cell[    1290] = 32'h2eef13e6;
    ram_cell[    1291] = 32'h15aa5fc7;
    ram_cell[    1292] = 32'h83d2e9aa;
    ram_cell[    1293] = 32'haa0c31ef;
    ram_cell[    1294] = 32'h2354b8c0;
    ram_cell[    1295] = 32'ha6eed6d0;
    ram_cell[    1296] = 32'hc9abffef;
    ram_cell[    1297] = 32'hd9d109c1;
    ram_cell[    1298] = 32'h7b01b86c;
    ram_cell[    1299] = 32'h18db87ff;
    ram_cell[    1300] = 32'h20acfcae;
    ram_cell[    1301] = 32'hd5a692e4;
    ram_cell[    1302] = 32'h103afce7;
    ram_cell[    1303] = 32'h700d09e0;
    ram_cell[    1304] = 32'h45196e43;
    ram_cell[    1305] = 32'h2e8cc53d;
    ram_cell[    1306] = 32'h9817e5bb;
    ram_cell[    1307] = 32'hf985cc4e;
    ram_cell[    1308] = 32'h3fc813a4;
    ram_cell[    1309] = 32'hea265b3a;
    ram_cell[    1310] = 32'h94440e05;
    ram_cell[    1311] = 32'h55327ba2;
    ram_cell[    1312] = 32'he239f400;
    ram_cell[    1313] = 32'hb7c65e0c;
    ram_cell[    1314] = 32'hfe4ce224;
    ram_cell[    1315] = 32'h7e68e51b;
    ram_cell[    1316] = 32'h03ad9890;
    ram_cell[    1317] = 32'h35cecdab;
    ram_cell[    1318] = 32'h1ca84346;
    ram_cell[    1319] = 32'h977d5ad4;
    ram_cell[    1320] = 32'hba685347;
    ram_cell[    1321] = 32'h6b175ac3;
    ram_cell[    1322] = 32'hfdb40b3e;
    ram_cell[    1323] = 32'h7b401a6f;
    ram_cell[    1324] = 32'h58a447aa;
    ram_cell[    1325] = 32'h92c6a587;
    ram_cell[    1326] = 32'h83c5ed41;
    ram_cell[    1327] = 32'hca5ee623;
    ram_cell[    1328] = 32'h9f939304;
    ram_cell[    1329] = 32'hf112d162;
    ram_cell[    1330] = 32'h540902c3;
    ram_cell[    1331] = 32'h352aab4f;
    ram_cell[    1332] = 32'hf2081108;
    ram_cell[    1333] = 32'hd18c07e2;
    ram_cell[    1334] = 32'h82262f49;
    ram_cell[    1335] = 32'h2232c806;
    ram_cell[    1336] = 32'ha3f90421;
    ram_cell[    1337] = 32'h02486bcb;
    ram_cell[    1338] = 32'h104c26c9;
    ram_cell[    1339] = 32'ha9bddf9d;
    ram_cell[    1340] = 32'h8a028bad;
    ram_cell[    1341] = 32'h9f852791;
    ram_cell[    1342] = 32'h8ee17c53;
    ram_cell[    1343] = 32'hbc852189;
    ram_cell[    1344] = 32'h671f9640;
    ram_cell[    1345] = 32'h49b1e23d;
    ram_cell[    1346] = 32'hf34f08e7;
    ram_cell[    1347] = 32'h01959f57;
    ram_cell[    1348] = 32'h3ff45354;
    ram_cell[    1349] = 32'h76511e2e;
    ram_cell[    1350] = 32'h85115440;
    ram_cell[    1351] = 32'h58bbceda;
    ram_cell[    1352] = 32'hfc97e2cf;
    ram_cell[    1353] = 32'h0eedc18b;
    ram_cell[    1354] = 32'hf65b8a51;
    ram_cell[    1355] = 32'h480477e3;
    ram_cell[    1356] = 32'he2bd29ea;
    ram_cell[    1357] = 32'hc48a6612;
    ram_cell[    1358] = 32'h6f0d01f5;
    ram_cell[    1359] = 32'hc9a38b61;
    ram_cell[    1360] = 32'hb6749e20;
    ram_cell[    1361] = 32'hdb56f038;
    ram_cell[    1362] = 32'hffdfb4cc;
    ram_cell[    1363] = 32'h32abdbd4;
    ram_cell[    1364] = 32'hce863e15;
    ram_cell[    1365] = 32'h60648c2c;
    ram_cell[    1366] = 32'hf7fe131c;
    ram_cell[    1367] = 32'he8f8e3c4;
    ram_cell[    1368] = 32'h98d0a6b7;
    ram_cell[    1369] = 32'h854c2e0e;
    ram_cell[    1370] = 32'h60154709;
    ram_cell[    1371] = 32'hd33667c0;
    ram_cell[    1372] = 32'h57199785;
    ram_cell[    1373] = 32'h9ae67067;
    ram_cell[    1374] = 32'hc2610fe7;
    ram_cell[    1375] = 32'h4e8cbda6;
    ram_cell[    1376] = 32'h71c087d8;
    ram_cell[    1377] = 32'h1f39a8bf;
    ram_cell[    1378] = 32'ha4fae3c3;
    ram_cell[    1379] = 32'hb1be587f;
    ram_cell[    1380] = 32'h864b8cf7;
    ram_cell[    1381] = 32'h56a8d5e1;
    ram_cell[    1382] = 32'h7e1106f2;
    ram_cell[    1383] = 32'h4f6f5ba4;
    ram_cell[    1384] = 32'h0cc26999;
    ram_cell[    1385] = 32'he20848b9;
    ram_cell[    1386] = 32'h3f87d07d;
    ram_cell[    1387] = 32'h22964c43;
    ram_cell[    1388] = 32'he0bd4775;
    ram_cell[    1389] = 32'h373fb2da;
    ram_cell[    1390] = 32'h3ca0dae6;
    ram_cell[    1391] = 32'hfdadffc0;
    ram_cell[    1392] = 32'h4def6c1a;
    ram_cell[    1393] = 32'h0885032f;
    ram_cell[    1394] = 32'h85998c7f;
    ram_cell[    1395] = 32'h531622cb;
    ram_cell[    1396] = 32'hd8014e0f;
    ram_cell[    1397] = 32'h467a7182;
    ram_cell[    1398] = 32'h064b59e1;
    ram_cell[    1399] = 32'he2b2b497;
    ram_cell[    1400] = 32'h1f5d87ee;
    ram_cell[    1401] = 32'h712479e9;
    ram_cell[    1402] = 32'h19b9195c;
    ram_cell[    1403] = 32'hca5da9e4;
    ram_cell[    1404] = 32'h3e46bc76;
    ram_cell[    1405] = 32'hee20ff78;
    ram_cell[    1406] = 32'hb9d94395;
    ram_cell[    1407] = 32'h87fa79ca;
    ram_cell[    1408] = 32'hd57bd1b0;
    ram_cell[    1409] = 32'h736417a2;
    ram_cell[    1410] = 32'hccfe4c5d;
    ram_cell[    1411] = 32'ha7fa9482;
    ram_cell[    1412] = 32'hd8bce75f;
    ram_cell[    1413] = 32'h892e991f;
    ram_cell[    1414] = 32'h2fb6dfb8;
    ram_cell[    1415] = 32'h5a093bd3;
    ram_cell[    1416] = 32'hc06fc5b8;
    ram_cell[    1417] = 32'h95293ae3;
    ram_cell[    1418] = 32'hf5025bf0;
    ram_cell[    1419] = 32'he6d4db61;
    ram_cell[    1420] = 32'h3cd35b56;
    ram_cell[    1421] = 32'h86b1e51d;
    ram_cell[    1422] = 32'h4a7a44c1;
    ram_cell[    1423] = 32'h899cccf3;
    ram_cell[    1424] = 32'h0d70c0e2;
    ram_cell[    1425] = 32'ha4519bec;
    ram_cell[    1426] = 32'hf07edaee;
    ram_cell[    1427] = 32'h3705db24;
    ram_cell[    1428] = 32'hd2a7cf5d;
    ram_cell[    1429] = 32'ha71a431d;
    ram_cell[    1430] = 32'ha604ed99;
    ram_cell[    1431] = 32'h875cb91d;
    ram_cell[    1432] = 32'h9f0f6b88;
    ram_cell[    1433] = 32'h7d3d495b;
    ram_cell[    1434] = 32'h06f4ace7;
    ram_cell[    1435] = 32'hdcf946da;
    ram_cell[    1436] = 32'hb0253752;
    ram_cell[    1437] = 32'haeae31fa;
    ram_cell[    1438] = 32'h7a509757;
    ram_cell[    1439] = 32'hed787982;
    ram_cell[    1440] = 32'ha14912ad;
    ram_cell[    1441] = 32'ha4e5f480;
    ram_cell[    1442] = 32'hcfa8a43c;
    ram_cell[    1443] = 32'h35a0e071;
    ram_cell[    1444] = 32'h5325f647;
    ram_cell[    1445] = 32'h95105672;
    ram_cell[    1446] = 32'h162b16f6;
    ram_cell[    1447] = 32'h4deeb07e;
    ram_cell[    1448] = 32'hed6b207a;
    ram_cell[    1449] = 32'hb4fe82d0;
    ram_cell[    1450] = 32'ha64c8406;
    ram_cell[    1451] = 32'hfd8c848c;
    ram_cell[    1452] = 32'h9f9c82df;
    ram_cell[    1453] = 32'h1ca6e91e;
    ram_cell[    1454] = 32'h819d8749;
    ram_cell[    1455] = 32'hfd0664d0;
    ram_cell[    1456] = 32'hccb229da;
    ram_cell[    1457] = 32'he0cae241;
    ram_cell[    1458] = 32'h9344004e;
    ram_cell[    1459] = 32'hbc8ddd55;
    ram_cell[    1460] = 32'haac084b3;
    ram_cell[    1461] = 32'ha2f4633f;
    ram_cell[    1462] = 32'hfa3b7068;
    ram_cell[    1463] = 32'h96fe202e;
    ram_cell[    1464] = 32'hf4fb952b;
    ram_cell[    1465] = 32'hf1ca0e1d;
    ram_cell[    1466] = 32'h6537d42c;
    ram_cell[    1467] = 32'h8b39e912;
    ram_cell[    1468] = 32'h7b1ffcb7;
    ram_cell[    1469] = 32'hb308ee33;
    ram_cell[    1470] = 32'h388cf3b3;
    ram_cell[    1471] = 32'hebdb6f36;
    ram_cell[    1472] = 32'ha87564df;
    ram_cell[    1473] = 32'ha2ec6280;
    ram_cell[    1474] = 32'h415cb039;
    ram_cell[    1475] = 32'h164a601a;
    ram_cell[    1476] = 32'hd55be0b4;
    ram_cell[    1477] = 32'hbdc4bc3b;
    ram_cell[    1478] = 32'h430eacd2;
    ram_cell[    1479] = 32'hdc77894b;
    ram_cell[    1480] = 32'h3eda62f6;
    ram_cell[    1481] = 32'ha5bccdc5;
    ram_cell[    1482] = 32'h070d3e4e;
    ram_cell[    1483] = 32'h21bccb7d;
    ram_cell[    1484] = 32'h3b37108f;
    ram_cell[    1485] = 32'h5a843bf9;
    ram_cell[    1486] = 32'h44b57a70;
    ram_cell[    1487] = 32'h4de8732b;
    ram_cell[    1488] = 32'h3c9421dd;
    ram_cell[    1489] = 32'hdec03395;
    ram_cell[    1490] = 32'hcef34d1d;
    ram_cell[    1491] = 32'heaaeaac8;
    ram_cell[    1492] = 32'hd6c7fdf2;
    ram_cell[    1493] = 32'h3e20cdf6;
    ram_cell[    1494] = 32'h26021cb1;
    ram_cell[    1495] = 32'h5603feb0;
    ram_cell[    1496] = 32'h1d52197e;
    ram_cell[    1497] = 32'h89e676a0;
    ram_cell[    1498] = 32'hc453b66d;
    ram_cell[    1499] = 32'h92454459;
    ram_cell[    1500] = 32'h75146922;
    ram_cell[    1501] = 32'h17a18fec;
    ram_cell[    1502] = 32'h90b4c691;
    ram_cell[    1503] = 32'hf9465cb3;
    ram_cell[    1504] = 32'he1cfdbec;
    ram_cell[    1505] = 32'hdb57ff90;
    ram_cell[    1506] = 32'h7490b035;
    ram_cell[    1507] = 32'hb3b4288e;
    ram_cell[    1508] = 32'h8330d603;
    ram_cell[    1509] = 32'hecbf4ccc;
    ram_cell[    1510] = 32'h08bc7fee;
    ram_cell[    1511] = 32'hf138161b;
    ram_cell[    1512] = 32'h62075dc2;
    ram_cell[    1513] = 32'ha9f77a6b;
    ram_cell[    1514] = 32'hb398f909;
    ram_cell[    1515] = 32'h807856cb;
    ram_cell[    1516] = 32'h228ea02f;
    ram_cell[    1517] = 32'hbc7946e1;
    ram_cell[    1518] = 32'h9da60ffe;
    ram_cell[    1519] = 32'h940c2825;
    ram_cell[    1520] = 32'h97035396;
    ram_cell[    1521] = 32'hbf71b5b1;
    ram_cell[    1522] = 32'h67d48bc8;
    ram_cell[    1523] = 32'h18bf5e7e;
    ram_cell[    1524] = 32'h223dd5c3;
    ram_cell[    1525] = 32'h710ba2ea;
    ram_cell[    1526] = 32'ha007b54a;
    ram_cell[    1527] = 32'hf6b20039;
    ram_cell[    1528] = 32'h415bb7d2;
    ram_cell[    1529] = 32'hb1f1a587;
    ram_cell[    1530] = 32'h3268b285;
    ram_cell[    1531] = 32'h18d18864;
    ram_cell[    1532] = 32'h6a7ca192;
    ram_cell[    1533] = 32'h2d124f8b;
    ram_cell[    1534] = 32'hfc2d1c1e;
    ram_cell[    1535] = 32'h6b030e90;
    ram_cell[    1536] = 32'h01b03211;
    ram_cell[    1537] = 32'hac3b98e0;
    ram_cell[    1538] = 32'h2ecc1113;
    ram_cell[    1539] = 32'hf8927ae5;
    ram_cell[    1540] = 32'h51e38add;
    ram_cell[    1541] = 32'ha74676b6;
    ram_cell[    1542] = 32'h1392b8e3;
    ram_cell[    1543] = 32'ha95b98a3;
    ram_cell[    1544] = 32'h6563139e;
    ram_cell[    1545] = 32'ha60213c5;
    ram_cell[    1546] = 32'h1b879c13;
    ram_cell[    1547] = 32'hf81c941c;
    ram_cell[    1548] = 32'h5a8f49f6;
    ram_cell[    1549] = 32'hbc3e8d69;
    ram_cell[    1550] = 32'h3b9ba81c;
    ram_cell[    1551] = 32'h7380b82f;
    ram_cell[    1552] = 32'h41039b5c;
    ram_cell[    1553] = 32'hbf0bad6c;
    ram_cell[    1554] = 32'h1cfc4b27;
    ram_cell[    1555] = 32'h5537ca74;
    ram_cell[    1556] = 32'h0537d61d;
    ram_cell[    1557] = 32'h16ddd238;
    ram_cell[    1558] = 32'h7c68303c;
    ram_cell[    1559] = 32'hd7c51e60;
    ram_cell[    1560] = 32'h19b195a3;
    ram_cell[    1561] = 32'h6f796191;
    ram_cell[    1562] = 32'h8adbc9bf;
    ram_cell[    1563] = 32'hd2b2e094;
    ram_cell[    1564] = 32'hd1a18c63;
    ram_cell[    1565] = 32'h47967cf1;
    ram_cell[    1566] = 32'h81b660a7;
    ram_cell[    1567] = 32'h746776e6;
    ram_cell[    1568] = 32'h25665edf;
    ram_cell[    1569] = 32'hd849acf7;
    ram_cell[    1570] = 32'h0c4c036b;
    ram_cell[    1571] = 32'h96d32dbb;
    ram_cell[    1572] = 32'h7ba7c139;
    ram_cell[    1573] = 32'hf74c90de;
    ram_cell[    1574] = 32'h0d6c319c;
    ram_cell[    1575] = 32'hb4bb0eb0;
    ram_cell[    1576] = 32'h78e7c282;
    ram_cell[    1577] = 32'h2f78d47b;
    ram_cell[    1578] = 32'h6867aa64;
    ram_cell[    1579] = 32'h04028cd5;
    ram_cell[    1580] = 32'h4ae5b6e1;
    ram_cell[    1581] = 32'hb86901d8;
    ram_cell[    1582] = 32'h2c1a2909;
    ram_cell[    1583] = 32'h5233ec5e;
    ram_cell[    1584] = 32'h818d6f0e;
    ram_cell[    1585] = 32'h4b34f7d5;
    ram_cell[    1586] = 32'ha20f0466;
    ram_cell[    1587] = 32'h3014b6ac;
    ram_cell[    1588] = 32'h6da8bedc;
    ram_cell[    1589] = 32'h123cbe7f;
    ram_cell[    1590] = 32'hcf93133e;
    ram_cell[    1591] = 32'h4e27df79;
    ram_cell[    1592] = 32'h83808cc4;
    ram_cell[    1593] = 32'h18c2baa7;
    ram_cell[    1594] = 32'h9d7fa53b;
    ram_cell[    1595] = 32'h744668d8;
    ram_cell[    1596] = 32'h02f9eea7;
    ram_cell[    1597] = 32'h2018cdfa;
    ram_cell[    1598] = 32'he2fda79a;
    ram_cell[    1599] = 32'hd4587dfd;
    ram_cell[    1600] = 32'h3c381422;
    ram_cell[    1601] = 32'hda87e2d5;
    ram_cell[    1602] = 32'h3f13a9c5;
    ram_cell[    1603] = 32'h764072a2;
    ram_cell[    1604] = 32'h1385d6fa;
    ram_cell[    1605] = 32'h8e29118d;
    ram_cell[    1606] = 32'h13f5e18f;
    ram_cell[    1607] = 32'ha9060b37;
    ram_cell[    1608] = 32'h6a6262af;
    ram_cell[    1609] = 32'h8953a4ac;
    ram_cell[    1610] = 32'h06be4fa7;
    ram_cell[    1611] = 32'h3e0ec17f;
    ram_cell[    1612] = 32'h4c1aca04;
    ram_cell[    1613] = 32'hccfcccbc;
    ram_cell[    1614] = 32'h4b9579ac;
    ram_cell[    1615] = 32'hfe421219;
    ram_cell[    1616] = 32'h4818f3a6;
    ram_cell[    1617] = 32'ha67a3ee9;
    ram_cell[    1618] = 32'he9064c3f;
    ram_cell[    1619] = 32'h84041bd3;
    ram_cell[    1620] = 32'h64df6b75;
    ram_cell[    1621] = 32'h7dd91788;
    ram_cell[    1622] = 32'h8f156f46;
    ram_cell[    1623] = 32'hc5a0b30c;
    ram_cell[    1624] = 32'h14dbb6df;
    ram_cell[    1625] = 32'hc6fb638a;
    ram_cell[    1626] = 32'hf2e624a6;
    ram_cell[    1627] = 32'hdaffc3a6;
    ram_cell[    1628] = 32'hee2fc26b;
    ram_cell[    1629] = 32'h260ca73e;
    ram_cell[    1630] = 32'h058667b1;
    ram_cell[    1631] = 32'h01d1c818;
    ram_cell[    1632] = 32'h0ff84f02;
    ram_cell[    1633] = 32'h99fae229;
    ram_cell[    1634] = 32'h99ac0bd0;
    ram_cell[    1635] = 32'hb0cae19a;
    ram_cell[    1636] = 32'hdc8465c4;
    ram_cell[    1637] = 32'h0b1fdf72;
    ram_cell[    1638] = 32'hfcc85c20;
    ram_cell[    1639] = 32'hc4186fbe;
    ram_cell[    1640] = 32'hc1eaaf93;
    ram_cell[    1641] = 32'h07710f67;
    ram_cell[    1642] = 32'h78a2d9a0;
    ram_cell[    1643] = 32'h4fc23ef2;
    ram_cell[    1644] = 32'hacc12e95;
    ram_cell[    1645] = 32'h1b3599be;
    ram_cell[    1646] = 32'h919d69a0;
    ram_cell[    1647] = 32'h4dd8ee74;
    ram_cell[    1648] = 32'hd011b460;
    ram_cell[    1649] = 32'h068bdf55;
    ram_cell[    1650] = 32'hc4596cdb;
    ram_cell[    1651] = 32'hc7bcfd88;
    ram_cell[    1652] = 32'hef347622;
    ram_cell[    1653] = 32'hf352d116;
    ram_cell[    1654] = 32'h8ce6a1c0;
    ram_cell[    1655] = 32'he8a602f5;
    ram_cell[    1656] = 32'h4460d0f8;
    ram_cell[    1657] = 32'hd7f6417b;
    ram_cell[    1658] = 32'h468b0641;
    ram_cell[    1659] = 32'habb1fc88;
    ram_cell[    1660] = 32'h214339a6;
    ram_cell[    1661] = 32'h95ffa888;
    ram_cell[    1662] = 32'h7fa21da3;
    ram_cell[    1663] = 32'h42560108;
    ram_cell[    1664] = 32'h9da0f135;
    ram_cell[    1665] = 32'h2050946f;
    ram_cell[    1666] = 32'h67cc5198;
    ram_cell[    1667] = 32'h9d755a24;
    ram_cell[    1668] = 32'hae5f9aca;
    ram_cell[    1669] = 32'h74d65e6d;
    ram_cell[    1670] = 32'hb8a73968;
    ram_cell[    1671] = 32'h20dcbe1d;
    ram_cell[    1672] = 32'h89347c10;
    ram_cell[    1673] = 32'h9dbbcfd8;
    ram_cell[    1674] = 32'hcd9ffbb5;
    ram_cell[    1675] = 32'hecae5be8;
    ram_cell[    1676] = 32'h91e557c9;
    ram_cell[    1677] = 32'h4719228b;
    ram_cell[    1678] = 32'h70c6439b;
    ram_cell[    1679] = 32'h9d21989a;
    ram_cell[    1680] = 32'h0d48d9a6;
    ram_cell[    1681] = 32'hf3356591;
    ram_cell[    1682] = 32'h6bf81fba;
    ram_cell[    1683] = 32'h1fde4c61;
    ram_cell[    1684] = 32'h93563682;
    ram_cell[    1685] = 32'h4f5fc3b3;
    ram_cell[    1686] = 32'hab42bb19;
    ram_cell[    1687] = 32'h22d78bc0;
    ram_cell[    1688] = 32'h69c4c33a;
    ram_cell[    1689] = 32'h6004f256;
    ram_cell[    1690] = 32'h3ddc8a46;
    ram_cell[    1691] = 32'hfa5e38c6;
    ram_cell[    1692] = 32'h56d4389d;
    ram_cell[    1693] = 32'h3adecfeb;
    ram_cell[    1694] = 32'h6c62932e;
    ram_cell[    1695] = 32'h2313bc26;
    ram_cell[    1696] = 32'h5852e1c6;
    ram_cell[    1697] = 32'h28086ae1;
    ram_cell[    1698] = 32'h68f99f97;
    ram_cell[    1699] = 32'h40589bb2;
    ram_cell[    1700] = 32'h8f3c7d92;
    ram_cell[    1701] = 32'hb8ca136a;
    ram_cell[    1702] = 32'h2aa4b986;
    ram_cell[    1703] = 32'h356275dd;
    ram_cell[    1704] = 32'h2cbc621e;
    ram_cell[    1705] = 32'h98be5557;
    ram_cell[    1706] = 32'h13e7b90f;
    ram_cell[    1707] = 32'h81152640;
    ram_cell[    1708] = 32'h53c5315f;
    ram_cell[    1709] = 32'h7287dd30;
    ram_cell[    1710] = 32'h77cfd5a8;
    ram_cell[    1711] = 32'hef0720a4;
    ram_cell[    1712] = 32'hb04b10f1;
    ram_cell[    1713] = 32'h6a99f402;
    ram_cell[    1714] = 32'h7a41c1d5;
    ram_cell[    1715] = 32'hf50fbcf4;
    ram_cell[    1716] = 32'h451074da;
    ram_cell[    1717] = 32'h63bdd05e;
    ram_cell[    1718] = 32'h599b4fe9;
    ram_cell[    1719] = 32'h4d747344;
    ram_cell[    1720] = 32'h705bb068;
    ram_cell[    1721] = 32'h80d9d2de;
    ram_cell[    1722] = 32'h677acbbe;
    ram_cell[    1723] = 32'h453aa3f8;
    ram_cell[    1724] = 32'h777efcd9;
    ram_cell[    1725] = 32'ha78ef18c;
    ram_cell[    1726] = 32'hd704b367;
    ram_cell[    1727] = 32'h1806d431;
    ram_cell[    1728] = 32'h565f85a6;
    ram_cell[    1729] = 32'h6d908f4f;
    ram_cell[    1730] = 32'h9a220a83;
    ram_cell[    1731] = 32'h3a29d93c;
    ram_cell[    1732] = 32'h6286b3fe;
    ram_cell[    1733] = 32'hb06e5aa2;
    ram_cell[    1734] = 32'ha21cafc4;
    ram_cell[    1735] = 32'h48d12c5f;
    ram_cell[    1736] = 32'h8553f63b;
    ram_cell[    1737] = 32'hdb4c0c36;
    ram_cell[    1738] = 32'h02e16f77;
    ram_cell[    1739] = 32'ha530133e;
    ram_cell[    1740] = 32'h07d4a00f;
    ram_cell[    1741] = 32'h4547f608;
    ram_cell[    1742] = 32'hb0c227d3;
    ram_cell[    1743] = 32'hacb394d4;
    ram_cell[    1744] = 32'h0a2f3157;
    ram_cell[    1745] = 32'heefa9cb1;
    ram_cell[    1746] = 32'hfc7f8506;
    ram_cell[    1747] = 32'h392fdc1c;
    ram_cell[    1748] = 32'hda117854;
    ram_cell[    1749] = 32'h76365652;
    ram_cell[    1750] = 32'h6fcf352b;
    ram_cell[    1751] = 32'h378b7e8e;
    ram_cell[    1752] = 32'hb8619e9c;
    ram_cell[    1753] = 32'h1bfbd5f0;
    ram_cell[    1754] = 32'h59a77e84;
    ram_cell[    1755] = 32'h7057aa6b;
    ram_cell[    1756] = 32'h2d14addd;
    ram_cell[    1757] = 32'ha80b125b;
    ram_cell[    1758] = 32'h130a9afb;
    ram_cell[    1759] = 32'hb50ee9ce;
    ram_cell[    1760] = 32'hf8ddf436;
    ram_cell[    1761] = 32'hea9773d6;
    ram_cell[    1762] = 32'h71058590;
    ram_cell[    1763] = 32'heca6f1bf;
    ram_cell[    1764] = 32'h9dac7a64;
    ram_cell[    1765] = 32'h6be9a918;
    ram_cell[    1766] = 32'h8126fecf;
    ram_cell[    1767] = 32'h9b6582da;
    ram_cell[    1768] = 32'hc485511c;
    ram_cell[    1769] = 32'h1e022f15;
    ram_cell[    1770] = 32'hc838d120;
    ram_cell[    1771] = 32'h6db2b100;
    ram_cell[    1772] = 32'h26129f38;
    ram_cell[    1773] = 32'h2395885d;
    ram_cell[    1774] = 32'hb8409b29;
    ram_cell[    1775] = 32'hd042d63f;
    ram_cell[    1776] = 32'hf9d9ef03;
    ram_cell[    1777] = 32'h04d23e9f;
    ram_cell[    1778] = 32'h0d0afd5d;
    ram_cell[    1779] = 32'h224a03ec;
    ram_cell[    1780] = 32'h0c424c18;
    ram_cell[    1781] = 32'hc093fa0d;
    ram_cell[    1782] = 32'h5310c2f6;
    ram_cell[    1783] = 32'he295765a;
    ram_cell[    1784] = 32'h7bebd8ed;
    ram_cell[    1785] = 32'hf4d7d914;
    ram_cell[    1786] = 32'h1497bdf8;
    ram_cell[    1787] = 32'h2029ba59;
    ram_cell[    1788] = 32'h705de62e;
    ram_cell[    1789] = 32'hc0923743;
    ram_cell[    1790] = 32'h6ad6187f;
    ram_cell[    1791] = 32'h65842e08;
    ram_cell[    1792] = 32'h9d0162a8;
    ram_cell[    1793] = 32'h56edebb1;
    ram_cell[    1794] = 32'h3cbda712;
    ram_cell[    1795] = 32'hbfb74cd0;
    ram_cell[    1796] = 32'h7a59717e;
    ram_cell[    1797] = 32'h724f3fc5;
    ram_cell[    1798] = 32'he77f8fa4;
    ram_cell[    1799] = 32'h73302410;
    ram_cell[    1800] = 32'h3d5436a9;
    ram_cell[    1801] = 32'h74240a2c;
    ram_cell[    1802] = 32'he2d9bd77;
    ram_cell[    1803] = 32'h92663ecd;
    ram_cell[    1804] = 32'h1a572d54;
    ram_cell[    1805] = 32'ha64df3e3;
    ram_cell[    1806] = 32'h7b79c2f5;
    ram_cell[    1807] = 32'hf6ee3edb;
    ram_cell[    1808] = 32'h4ac81e89;
    ram_cell[    1809] = 32'h8d1dc424;
    ram_cell[    1810] = 32'ha90fb1c8;
    ram_cell[    1811] = 32'h835f7920;
    ram_cell[    1812] = 32'he72e880d;
    ram_cell[    1813] = 32'hccabec82;
    ram_cell[    1814] = 32'h2e71edea;
    ram_cell[    1815] = 32'h840e7c1c;
    ram_cell[    1816] = 32'hf03aa91f;
    ram_cell[    1817] = 32'h1bdb973f;
    ram_cell[    1818] = 32'hc8070ba7;
    ram_cell[    1819] = 32'hf4fbba8b;
    ram_cell[    1820] = 32'h46ee7254;
    ram_cell[    1821] = 32'hd2add3e8;
    ram_cell[    1822] = 32'h140b1dbc;
    ram_cell[    1823] = 32'h26553e13;
    ram_cell[    1824] = 32'h601a5d58;
    ram_cell[    1825] = 32'hab0ea3cc;
    ram_cell[    1826] = 32'h5ff432b7;
    ram_cell[    1827] = 32'ha6062680;
    ram_cell[    1828] = 32'hfc92989d;
    ram_cell[    1829] = 32'h2aedf03a;
    ram_cell[    1830] = 32'h2d1a1016;
    ram_cell[    1831] = 32'he8baf50a;
    ram_cell[    1832] = 32'h4c8bd9b3;
    ram_cell[    1833] = 32'h44a3c5c5;
    ram_cell[    1834] = 32'h07f31842;
    ram_cell[    1835] = 32'h48c9f023;
    ram_cell[    1836] = 32'hc25e19fc;
    ram_cell[    1837] = 32'h61964881;
    ram_cell[    1838] = 32'hca680645;
    ram_cell[    1839] = 32'hfd8d5390;
    ram_cell[    1840] = 32'h880b2282;
    ram_cell[    1841] = 32'hb463e880;
    ram_cell[    1842] = 32'hcd849467;
    ram_cell[    1843] = 32'haf54ec14;
    ram_cell[    1844] = 32'h1b28c619;
    ram_cell[    1845] = 32'h6eef6b5d;
    ram_cell[    1846] = 32'h08755def;
    ram_cell[    1847] = 32'h2103aaaa;
    ram_cell[    1848] = 32'h9f9c8c24;
    ram_cell[    1849] = 32'hc9bd63e9;
    ram_cell[    1850] = 32'h5dbc1e84;
    ram_cell[    1851] = 32'hef49e8b9;
    ram_cell[    1852] = 32'h09604d02;
    ram_cell[    1853] = 32'h249002a1;
    ram_cell[    1854] = 32'haff15567;
    ram_cell[    1855] = 32'h767dc76f;
    ram_cell[    1856] = 32'ha5b222aa;
    ram_cell[    1857] = 32'h60ffcf4e;
    ram_cell[    1858] = 32'hfddfbc50;
    ram_cell[    1859] = 32'h1cadcfe3;
    ram_cell[    1860] = 32'h48421aa1;
    ram_cell[    1861] = 32'hf011dd68;
    ram_cell[    1862] = 32'hacc4e183;
    ram_cell[    1863] = 32'h92d8d8fa;
    ram_cell[    1864] = 32'h9fbc5592;
    ram_cell[    1865] = 32'h25063795;
    ram_cell[    1866] = 32'hfe80923e;
    ram_cell[    1867] = 32'habcbfdef;
    ram_cell[    1868] = 32'h9fdd3afa;
    ram_cell[    1869] = 32'h369d0305;
    ram_cell[    1870] = 32'h9227e3df;
    ram_cell[    1871] = 32'hcbff07b2;
    ram_cell[    1872] = 32'h513b66d8;
    ram_cell[    1873] = 32'h450962c6;
    ram_cell[    1874] = 32'h5e42d8df;
    ram_cell[    1875] = 32'he975823d;
    ram_cell[    1876] = 32'h7aa24f7d;
    ram_cell[    1877] = 32'h5634b0fa;
    ram_cell[    1878] = 32'ha18e15c4;
    ram_cell[    1879] = 32'hb0526d88;
    ram_cell[    1880] = 32'h049acf8d;
    ram_cell[    1881] = 32'hedf4575a;
    ram_cell[    1882] = 32'h13b187c7;
    ram_cell[    1883] = 32'h4546312b;
    ram_cell[    1884] = 32'h3ed14175;
    ram_cell[    1885] = 32'hce56cc70;
    ram_cell[    1886] = 32'hbf4c4d0b;
    ram_cell[    1887] = 32'h74b98483;
    ram_cell[    1888] = 32'ha0a4bbbe;
    ram_cell[    1889] = 32'h2c594af4;
    ram_cell[    1890] = 32'h6cc2934d;
    ram_cell[    1891] = 32'hb961cf21;
    ram_cell[    1892] = 32'h475eafbd;
    ram_cell[    1893] = 32'h4b68c5de;
    ram_cell[    1894] = 32'hd5a8a653;
    ram_cell[    1895] = 32'hd5bdf669;
    ram_cell[    1896] = 32'hfde26e0f;
    ram_cell[    1897] = 32'hf4ad5a50;
    ram_cell[    1898] = 32'h080764c7;
    ram_cell[    1899] = 32'hcf46d79d;
    ram_cell[    1900] = 32'hcb2288f4;
    ram_cell[    1901] = 32'h12bc7970;
    ram_cell[    1902] = 32'hab7916b6;
    ram_cell[    1903] = 32'h609a6a9c;
    ram_cell[    1904] = 32'h679d2c1f;
    ram_cell[    1905] = 32'he2403b6f;
    ram_cell[    1906] = 32'h4761fea5;
    ram_cell[    1907] = 32'h56061d87;
    ram_cell[    1908] = 32'habde6bc5;
    ram_cell[    1909] = 32'hd4bdf6e2;
    ram_cell[    1910] = 32'hf90e8f5b;
    ram_cell[    1911] = 32'h8bafa989;
    ram_cell[    1912] = 32'h678be15d;
    ram_cell[    1913] = 32'h60338aac;
    ram_cell[    1914] = 32'h55540ac1;
    ram_cell[    1915] = 32'h4b7f26bc;
    ram_cell[    1916] = 32'h62c5f26c;
    ram_cell[    1917] = 32'h18ce2555;
    ram_cell[    1918] = 32'h984b86e9;
    ram_cell[    1919] = 32'h002b175f;
    ram_cell[    1920] = 32'ha623f841;
    ram_cell[    1921] = 32'h13dc3e39;
    ram_cell[    1922] = 32'ha2a0d434;
    ram_cell[    1923] = 32'hb373fc06;
    ram_cell[    1924] = 32'h217c3e50;
    ram_cell[    1925] = 32'hab484740;
    ram_cell[    1926] = 32'h8f971527;
    ram_cell[    1927] = 32'h2a07321c;
    ram_cell[    1928] = 32'ha0dc6877;
    ram_cell[    1929] = 32'h233db323;
    ram_cell[    1930] = 32'h6b152307;
    ram_cell[    1931] = 32'h2e987798;
    ram_cell[    1932] = 32'he5e04537;
    ram_cell[    1933] = 32'h5a3e9802;
    ram_cell[    1934] = 32'hc7be17f5;
    ram_cell[    1935] = 32'h5ba0dac2;
    ram_cell[    1936] = 32'hf4a658a4;
    ram_cell[    1937] = 32'had25d241;
    ram_cell[    1938] = 32'hbff158c8;
    ram_cell[    1939] = 32'he77cc7a9;
    ram_cell[    1940] = 32'h78f98990;
    ram_cell[    1941] = 32'h626b1d98;
    ram_cell[    1942] = 32'h1390720b;
    ram_cell[    1943] = 32'h1f32dd52;
    ram_cell[    1944] = 32'ha5392ddb;
    ram_cell[    1945] = 32'h0b8b8b71;
    ram_cell[    1946] = 32'had7fe13f;
    ram_cell[    1947] = 32'h9897f629;
    ram_cell[    1948] = 32'h1670623f;
    ram_cell[    1949] = 32'h01b689b1;
    ram_cell[    1950] = 32'h6c082b38;
    ram_cell[    1951] = 32'h6021e5d8;
    ram_cell[    1952] = 32'hef4c6284;
    ram_cell[    1953] = 32'hc373b70f;
    ram_cell[    1954] = 32'h7ea453de;
    ram_cell[    1955] = 32'h562dcac0;
    ram_cell[    1956] = 32'ha76a7af8;
    ram_cell[    1957] = 32'h0c0c3f85;
    ram_cell[    1958] = 32'h23e336cd;
    ram_cell[    1959] = 32'ha6ec997e;
    ram_cell[    1960] = 32'he0e7a12d;
    ram_cell[    1961] = 32'haf0effa3;
    ram_cell[    1962] = 32'hfdb9aec7;
    ram_cell[    1963] = 32'hd00efb22;
    ram_cell[    1964] = 32'h9e26c729;
    ram_cell[    1965] = 32'h4d909154;
    ram_cell[    1966] = 32'hb171a1c0;
    ram_cell[    1967] = 32'h5199227d;
    ram_cell[    1968] = 32'hb617d8a8;
    ram_cell[    1969] = 32'h8cb107d8;
    ram_cell[    1970] = 32'hacec6b61;
    ram_cell[    1971] = 32'hbb0b4b61;
    ram_cell[    1972] = 32'hef6f7a3a;
    ram_cell[    1973] = 32'h9dcc13d4;
    ram_cell[    1974] = 32'hc445e491;
    ram_cell[    1975] = 32'h2a7a555a;
    ram_cell[    1976] = 32'hacc016ce;
    ram_cell[    1977] = 32'h464523c6;
    ram_cell[    1978] = 32'h877d087d;
    ram_cell[    1979] = 32'hce8b76f9;
    ram_cell[    1980] = 32'h3483f2fb;
    ram_cell[    1981] = 32'hf8329243;
    ram_cell[    1982] = 32'h6f9f0b15;
    ram_cell[    1983] = 32'h2f9d7175;
    ram_cell[    1984] = 32'h7a5aa8aa;
    ram_cell[    1985] = 32'h0acded40;
    ram_cell[    1986] = 32'hf60c0ced;
    ram_cell[    1987] = 32'h81b716b9;
    ram_cell[    1988] = 32'h0bcf4ecf;
    ram_cell[    1989] = 32'hf5bf3e34;
    ram_cell[    1990] = 32'h0e505ffe;
    ram_cell[    1991] = 32'ha3fe6576;
    ram_cell[    1992] = 32'h416beabe;
    ram_cell[    1993] = 32'hb2e09dfb;
    ram_cell[    1994] = 32'h7e6b7928;
    ram_cell[    1995] = 32'h97541a3f;
    ram_cell[    1996] = 32'hea229d6d;
    ram_cell[    1997] = 32'h04b74a37;
    ram_cell[    1998] = 32'h18a0f788;
    ram_cell[    1999] = 32'h1eb115ef;
    ram_cell[    2000] = 32'h5cc5ad8f;
    ram_cell[    2001] = 32'heb3156bb;
    ram_cell[    2002] = 32'h149955c5;
    ram_cell[    2003] = 32'h4ba94356;
    ram_cell[    2004] = 32'h1f403644;
    ram_cell[    2005] = 32'h25e4bd8c;
    ram_cell[    2006] = 32'hbbbe84b6;
    ram_cell[    2007] = 32'hc9eab787;
    ram_cell[    2008] = 32'h92123bfe;
    ram_cell[    2009] = 32'h4449d5b2;
    ram_cell[    2010] = 32'h407496aa;
    ram_cell[    2011] = 32'h91451e3a;
    ram_cell[    2012] = 32'h0920562d;
    ram_cell[    2013] = 32'h9d5d9e6d;
    ram_cell[    2014] = 32'hb5626961;
    ram_cell[    2015] = 32'hb56be083;
    ram_cell[    2016] = 32'hab3ecf4f;
    ram_cell[    2017] = 32'h9dd39b6b;
    ram_cell[    2018] = 32'h34a8f65f;
    ram_cell[    2019] = 32'he9530ce7;
    ram_cell[    2020] = 32'hd671a83c;
    ram_cell[    2021] = 32'h17e85981;
    ram_cell[    2022] = 32'h4279da9a;
    ram_cell[    2023] = 32'ha7efd18b;
    ram_cell[    2024] = 32'hf89a4c28;
    ram_cell[    2025] = 32'h1b8bf4f2;
    ram_cell[    2026] = 32'h2394f9d6;
    ram_cell[    2027] = 32'h43cb8fd3;
    ram_cell[    2028] = 32'h70e6a119;
    ram_cell[    2029] = 32'h54f1d1bc;
    ram_cell[    2030] = 32'hfbc979f5;
    ram_cell[    2031] = 32'h8266f8ab;
    ram_cell[    2032] = 32'h19ccba83;
    ram_cell[    2033] = 32'ha9e7d007;
    ram_cell[    2034] = 32'hffb3f2c6;
    ram_cell[    2035] = 32'h376d41bc;
    ram_cell[    2036] = 32'hb1066e58;
    ram_cell[    2037] = 32'h36c98bc8;
    ram_cell[    2038] = 32'h92ad0088;
    ram_cell[    2039] = 32'h5573ee21;
    ram_cell[    2040] = 32'h77f59238;
    ram_cell[    2041] = 32'h4fdef196;
    ram_cell[    2042] = 32'h1ed951e2;
    ram_cell[    2043] = 32'h6801c18a;
    ram_cell[    2044] = 32'h184763db;
    ram_cell[    2045] = 32'h68ded6d5;
    ram_cell[    2046] = 32'h27dc6ef4;
    ram_cell[    2047] = 32'h1f75edd8;
    // src matrix B
    ram_cell[    2048] = 32'h0c6802fa;
    ram_cell[    2049] = 32'h87140949;
    ram_cell[    2050] = 32'hb3621657;
    ram_cell[    2051] = 32'haddfc230;
    ram_cell[    2052] = 32'h969b2d8a;
    ram_cell[    2053] = 32'hc922f615;
    ram_cell[    2054] = 32'h331d71b4;
    ram_cell[    2055] = 32'h7cdc9659;
    ram_cell[    2056] = 32'h9b522a4a;
    ram_cell[    2057] = 32'h3995f6b4;
    ram_cell[    2058] = 32'h812b718e;
    ram_cell[    2059] = 32'hc5d81ccf;
    ram_cell[    2060] = 32'he890f2cc;
    ram_cell[    2061] = 32'h910148f3;
    ram_cell[    2062] = 32'h418e6583;
    ram_cell[    2063] = 32'hc84128c5;
    ram_cell[    2064] = 32'h433080e2;
    ram_cell[    2065] = 32'h25c4c58b;
    ram_cell[    2066] = 32'hef294dca;
    ram_cell[    2067] = 32'hcc6beec0;
    ram_cell[    2068] = 32'h574db0c4;
    ram_cell[    2069] = 32'hb2c73bb5;
    ram_cell[    2070] = 32'hb07799a7;
    ram_cell[    2071] = 32'h8dd1b046;
    ram_cell[    2072] = 32'h15b0e67e;
    ram_cell[    2073] = 32'h2f5feacb;
    ram_cell[    2074] = 32'h584284b4;
    ram_cell[    2075] = 32'h41f0dd13;
    ram_cell[    2076] = 32'h962d2ef3;
    ram_cell[    2077] = 32'hf856c8d2;
    ram_cell[    2078] = 32'h2f740607;
    ram_cell[    2079] = 32'h29dc36c1;
    ram_cell[    2080] = 32'hc84d005e;
    ram_cell[    2081] = 32'h2b4c0ceb;
    ram_cell[    2082] = 32'h68ba37bf;
    ram_cell[    2083] = 32'h2015a961;
    ram_cell[    2084] = 32'h0be790fc;
    ram_cell[    2085] = 32'haa72275d;
    ram_cell[    2086] = 32'h7a2d19a5;
    ram_cell[    2087] = 32'h6b7b597f;
    ram_cell[    2088] = 32'he6f771a7;
    ram_cell[    2089] = 32'h9af17fdf;
    ram_cell[    2090] = 32'h5e4c6a79;
    ram_cell[    2091] = 32'hb5426a41;
    ram_cell[    2092] = 32'h064d8734;
    ram_cell[    2093] = 32'h8a8a67b4;
    ram_cell[    2094] = 32'h0d137d6a;
    ram_cell[    2095] = 32'h04ab51d4;
    ram_cell[    2096] = 32'hc8cf59e7;
    ram_cell[    2097] = 32'hfdeb4cbe;
    ram_cell[    2098] = 32'h272afe5e;
    ram_cell[    2099] = 32'h8b187cb2;
    ram_cell[    2100] = 32'hf0b065c6;
    ram_cell[    2101] = 32'h165c5283;
    ram_cell[    2102] = 32'hbb457615;
    ram_cell[    2103] = 32'h0d7ab225;
    ram_cell[    2104] = 32'hfaf531ee;
    ram_cell[    2105] = 32'haca76e7c;
    ram_cell[    2106] = 32'h93202ea5;
    ram_cell[    2107] = 32'h4883487e;
    ram_cell[    2108] = 32'h94f5be6c;
    ram_cell[    2109] = 32'h68277ccb;
    ram_cell[    2110] = 32'hf003aec8;
    ram_cell[    2111] = 32'h042b7230;
    ram_cell[    2112] = 32'hddb7fd94;
    ram_cell[    2113] = 32'h4e797145;
    ram_cell[    2114] = 32'h4bd2a519;
    ram_cell[    2115] = 32'h17ac48f1;
    ram_cell[    2116] = 32'hee70a64d;
    ram_cell[    2117] = 32'h48a0ca48;
    ram_cell[    2118] = 32'h34654cf1;
    ram_cell[    2119] = 32'h0904748d;
    ram_cell[    2120] = 32'h9c40af94;
    ram_cell[    2121] = 32'hdd9cab15;
    ram_cell[    2122] = 32'hb3f90c7e;
    ram_cell[    2123] = 32'h0892ed75;
    ram_cell[    2124] = 32'h94b25530;
    ram_cell[    2125] = 32'hb16c0e8d;
    ram_cell[    2126] = 32'he4347924;
    ram_cell[    2127] = 32'h54737524;
    ram_cell[    2128] = 32'h065a79b6;
    ram_cell[    2129] = 32'h87b50b8d;
    ram_cell[    2130] = 32'h932d32fe;
    ram_cell[    2131] = 32'haab3265b;
    ram_cell[    2132] = 32'h09b1f537;
    ram_cell[    2133] = 32'hcc38405b;
    ram_cell[    2134] = 32'h59f2aad6;
    ram_cell[    2135] = 32'h5685f644;
    ram_cell[    2136] = 32'ha32f7de0;
    ram_cell[    2137] = 32'hfa64926e;
    ram_cell[    2138] = 32'hcd6a0219;
    ram_cell[    2139] = 32'h861f1f98;
    ram_cell[    2140] = 32'hfba89686;
    ram_cell[    2141] = 32'h442312f0;
    ram_cell[    2142] = 32'h0a42518e;
    ram_cell[    2143] = 32'hc17f4128;
    ram_cell[    2144] = 32'h3fa6c326;
    ram_cell[    2145] = 32'hdf42e0ce;
    ram_cell[    2146] = 32'h8e78fdd4;
    ram_cell[    2147] = 32'hc54abe8e;
    ram_cell[    2148] = 32'h708ddb86;
    ram_cell[    2149] = 32'he1636b06;
    ram_cell[    2150] = 32'h6d50477b;
    ram_cell[    2151] = 32'hafe36ceb;
    ram_cell[    2152] = 32'h9a4efde2;
    ram_cell[    2153] = 32'h3be16f6a;
    ram_cell[    2154] = 32'h0237d2ad;
    ram_cell[    2155] = 32'hd0d252b0;
    ram_cell[    2156] = 32'h5ff66323;
    ram_cell[    2157] = 32'h7768924a;
    ram_cell[    2158] = 32'hd98205ba;
    ram_cell[    2159] = 32'heb985f4a;
    ram_cell[    2160] = 32'h1ae44af9;
    ram_cell[    2161] = 32'hdd1ea688;
    ram_cell[    2162] = 32'hfcafa0aa;
    ram_cell[    2163] = 32'h1ea086ba;
    ram_cell[    2164] = 32'h0b225cf4;
    ram_cell[    2165] = 32'hcc69c6b4;
    ram_cell[    2166] = 32'hb35ba602;
    ram_cell[    2167] = 32'h8e6600e0;
    ram_cell[    2168] = 32'hcb712ae5;
    ram_cell[    2169] = 32'hb44b3159;
    ram_cell[    2170] = 32'h60a70db3;
    ram_cell[    2171] = 32'hf3d3ad51;
    ram_cell[    2172] = 32'hd54f7b49;
    ram_cell[    2173] = 32'h9e851955;
    ram_cell[    2174] = 32'hea5af2cb;
    ram_cell[    2175] = 32'h5eb215dd;
    ram_cell[    2176] = 32'hc3241edb;
    ram_cell[    2177] = 32'hc0a3d53e;
    ram_cell[    2178] = 32'h702dca62;
    ram_cell[    2179] = 32'h47b5f9da;
    ram_cell[    2180] = 32'h685ec292;
    ram_cell[    2181] = 32'h37c8aa28;
    ram_cell[    2182] = 32'he4f81f3e;
    ram_cell[    2183] = 32'ha1de1604;
    ram_cell[    2184] = 32'h97265561;
    ram_cell[    2185] = 32'h6ad0b2e4;
    ram_cell[    2186] = 32'hfbbaa352;
    ram_cell[    2187] = 32'hdd6b635d;
    ram_cell[    2188] = 32'h18eef9d4;
    ram_cell[    2189] = 32'hc71a4674;
    ram_cell[    2190] = 32'hfac70337;
    ram_cell[    2191] = 32'h5324a117;
    ram_cell[    2192] = 32'hbfe9cd74;
    ram_cell[    2193] = 32'h8350238d;
    ram_cell[    2194] = 32'h8e0cad96;
    ram_cell[    2195] = 32'hd0c5f84f;
    ram_cell[    2196] = 32'h83f03412;
    ram_cell[    2197] = 32'h94b4a1d9;
    ram_cell[    2198] = 32'hc733b5f1;
    ram_cell[    2199] = 32'h2d889a1b;
    ram_cell[    2200] = 32'h30351f61;
    ram_cell[    2201] = 32'he10d884f;
    ram_cell[    2202] = 32'hb4e6c0b1;
    ram_cell[    2203] = 32'he2cd12fe;
    ram_cell[    2204] = 32'h443edbb6;
    ram_cell[    2205] = 32'he5663739;
    ram_cell[    2206] = 32'hce96547a;
    ram_cell[    2207] = 32'hffb30a2c;
    ram_cell[    2208] = 32'h0f9da53c;
    ram_cell[    2209] = 32'h954fd0ac;
    ram_cell[    2210] = 32'h5d15a99f;
    ram_cell[    2211] = 32'h4ea30d04;
    ram_cell[    2212] = 32'hc9ab4c9b;
    ram_cell[    2213] = 32'hb883f3cc;
    ram_cell[    2214] = 32'hc3526cdc;
    ram_cell[    2215] = 32'ha874f4cb;
    ram_cell[    2216] = 32'h84ed7bba;
    ram_cell[    2217] = 32'h93df5bda;
    ram_cell[    2218] = 32'h1dd6c748;
    ram_cell[    2219] = 32'h1d8f99f6;
    ram_cell[    2220] = 32'h2d256d2f;
    ram_cell[    2221] = 32'h02705b5e;
    ram_cell[    2222] = 32'h1a90dbf2;
    ram_cell[    2223] = 32'hc223a825;
    ram_cell[    2224] = 32'h7212335a;
    ram_cell[    2225] = 32'h651dfc04;
    ram_cell[    2226] = 32'h67e6bce2;
    ram_cell[    2227] = 32'he6b2edfd;
    ram_cell[    2228] = 32'hfdf38445;
    ram_cell[    2229] = 32'hf7cf3ccc;
    ram_cell[    2230] = 32'had82990c;
    ram_cell[    2231] = 32'hc00cb9f7;
    ram_cell[    2232] = 32'hdcbf4595;
    ram_cell[    2233] = 32'h6fc835b5;
    ram_cell[    2234] = 32'h003761c4;
    ram_cell[    2235] = 32'h12795077;
    ram_cell[    2236] = 32'h41feff60;
    ram_cell[    2237] = 32'h3a6da7c5;
    ram_cell[    2238] = 32'hf57942ee;
    ram_cell[    2239] = 32'h779b0bfc;
    ram_cell[    2240] = 32'hd09601a6;
    ram_cell[    2241] = 32'h695a91f7;
    ram_cell[    2242] = 32'hf28887b4;
    ram_cell[    2243] = 32'h43a5ded2;
    ram_cell[    2244] = 32'h6334bc3a;
    ram_cell[    2245] = 32'hc13ee686;
    ram_cell[    2246] = 32'hc1d1b95a;
    ram_cell[    2247] = 32'h60708eeb;
    ram_cell[    2248] = 32'hb3274ed2;
    ram_cell[    2249] = 32'h2eec45a3;
    ram_cell[    2250] = 32'h861fb071;
    ram_cell[    2251] = 32'h6753dee2;
    ram_cell[    2252] = 32'h0aa42c98;
    ram_cell[    2253] = 32'h2e439f9b;
    ram_cell[    2254] = 32'h9597e9ef;
    ram_cell[    2255] = 32'hefa8385c;
    ram_cell[    2256] = 32'h3a92754c;
    ram_cell[    2257] = 32'h4b1f68fe;
    ram_cell[    2258] = 32'h9e395b06;
    ram_cell[    2259] = 32'haa05767c;
    ram_cell[    2260] = 32'h29002ff4;
    ram_cell[    2261] = 32'hae4fabe5;
    ram_cell[    2262] = 32'hb4c3e7e2;
    ram_cell[    2263] = 32'ha0155296;
    ram_cell[    2264] = 32'h3b142782;
    ram_cell[    2265] = 32'h835dfd07;
    ram_cell[    2266] = 32'h1a8725c3;
    ram_cell[    2267] = 32'hce95b1d6;
    ram_cell[    2268] = 32'h7dadc64e;
    ram_cell[    2269] = 32'h682cec43;
    ram_cell[    2270] = 32'ha14cfd2e;
    ram_cell[    2271] = 32'hbc6beb2c;
    ram_cell[    2272] = 32'he3174d43;
    ram_cell[    2273] = 32'h4ecac114;
    ram_cell[    2274] = 32'h6147c872;
    ram_cell[    2275] = 32'haa8f85f4;
    ram_cell[    2276] = 32'h6a66462d;
    ram_cell[    2277] = 32'h1e3a6b8d;
    ram_cell[    2278] = 32'h5307594a;
    ram_cell[    2279] = 32'h3bedf3ff;
    ram_cell[    2280] = 32'hc2393c59;
    ram_cell[    2281] = 32'h2c2ad2ce;
    ram_cell[    2282] = 32'h3b19158e;
    ram_cell[    2283] = 32'hb6132805;
    ram_cell[    2284] = 32'hdd8b4277;
    ram_cell[    2285] = 32'h9647c30a;
    ram_cell[    2286] = 32'h4a0b0163;
    ram_cell[    2287] = 32'hf41ac517;
    ram_cell[    2288] = 32'hc5c09a6a;
    ram_cell[    2289] = 32'he0dfc914;
    ram_cell[    2290] = 32'h7bbaab50;
    ram_cell[    2291] = 32'h7827afb8;
    ram_cell[    2292] = 32'hd32cbbea;
    ram_cell[    2293] = 32'heb056405;
    ram_cell[    2294] = 32'h476b3ca5;
    ram_cell[    2295] = 32'h8a222b68;
    ram_cell[    2296] = 32'h08fcb451;
    ram_cell[    2297] = 32'hab03daf9;
    ram_cell[    2298] = 32'h230589db;
    ram_cell[    2299] = 32'hcc9f32c9;
    ram_cell[    2300] = 32'h44500e52;
    ram_cell[    2301] = 32'ha23a3280;
    ram_cell[    2302] = 32'h9cef1f4b;
    ram_cell[    2303] = 32'h30cd2feb;
    ram_cell[    2304] = 32'h729b063c;
    ram_cell[    2305] = 32'h8a26e234;
    ram_cell[    2306] = 32'h7708d89c;
    ram_cell[    2307] = 32'hfebf1bf2;
    ram_cell[    2308] = 32'h21cda2a3;
    ram_cell[    2309] = 32'h57adebff;
    ram_cell[    2310] = 32'h1690d3ec;
    ram_cell[    2311] = 32'hf7ad82ad;
    ram_cell[    2312] = 32'h6c460f7b;
    ram_cell[    2313] = 32'he704000e;
    ram_cell[    2314] = 32'h5d890080;
    ram_cell[    2315] = 32'hb0bfdeeb;
    ram_cell[    2316] = 32'hc08e6ab0;
    ram_cell[    2317] = 32'h58457d76;
    ram_cell[    2318] = 32'h633f94f7;
    ram_cell[    2319] = 32'hdc9e1f5a;
    ram_cell[    2320] = 32'h3ddd1879;
    ram_cell[    2321] = 32'h4ae8c0a4;
    ram_cell[    2322] = 32'h6baa162c;
    ram_cell[    2323] = 32'h0275195a;
    ram_cell[    2324] = 32'h526ece53;
    ram_cell[    2325] = 32'h7cf74cec;
    ram_cell[    2326] = 32'h3e92601b;
    ram_cell[    2327] = 32'hc2d5e4a4;
    ram_cell[    2328] = 32'h562219eb;
    ram_cell[    2329] = 32'h35d98157;
    ram_cell[    2330] = 32'hcdf57591;
    ram_cell[    2331] = 32'h52e66f84;
    ram_cell[    2332] = 32'hc054231d;
    ram_cell[    2333] = 32'h6622c342;
    ram_cell[    2334] = 32'hd1f738ac;
    ram_cell[    2335] = 32'hf04fd2f3;
    ram_cell[    2336] = 32'h51a8d6ec;
    ram_cell[    2337] = 32'hac6f7470;
    ram_cell[    2338] = 32'h3106dff1;
    ram_cell[    2339] = 32'he28dc81b;
    ram_cell[    2340] = 32'h87566b42;
    ram_cell[    2341] = 32'h75534acf;
    ram_cell[    2342] = 32'h42a6e3f0;
    ram_cell[    2343] = 32'h5fd737c6;
    ram_cell[    2344] = 32'hcac35ceb;
    ram_cell[    2345] = 32'h3105fad5;
    ram_cell[    2346] = 32'h5eb1ca25;
    ram_cell[    2347] = 32'h57454fef;
    ram_cell[    2348] = 32'h1350d03f;
    ram_cell[    2349] = 32'h54f32be5;
    ram_cell[    2350] = 32'hd2c02d2e;
    ram_cell[    2351] = 32'h9e4c00b8;
    ram_cell[    2352] = 32'hfce585cf;
    ram_cell[    2353] = 32'h3522f074;
    ram_cell[    2354] = 32'hdad544e0;
    ram_cell[    2355] = 32'h33f93c23;
    ram_cell[    2356] = 32'hcae96bdd;
    ram_cell[    2357] = 32'hbf15546e;
    ram_cell[    2358] = 32'h3b4c0ced;
    ram_cell[    2359] = 32'h42d43c0a;
    ram_cell[    2360] = 32'h414a7cec;
    ram_cell[    2361] = 32'hfda73bca;
    ram_cell[    2362] = 32'ha6998eac;
    ram_cell[    2363] = 32'h318683c9;
    ram_cell[    2364] = 32'h699bcbbf;
    ram_cell[    2365] = 32'h80fe0891;
    ram_cell[    2366] = 32'he3b76c69;
    ram_cell[    2367] = 32'h9a272def;
    ram_cell[    2368] = 32'h39cd5bfe;
    ram_cell[    2369] = 32'h97675813;
    ram_cell[    2370] = 32'h396504e0;
    ram_cell[    2371] = 32'he19f9c61;
    ram_cell[    2372] = 32'h44f9dec6;
    ram_cell[    2373] = 32'h40f97551;
    ram_cell[    2374] = 32'h0db1e516;
    ram_cell[    2375] = 32'h23124ca0;
    ram_cell[    2376] = 32'h92defb69;
    ram_cell[    2377] = 32'h9b64979c;
    ram_cell[    2378] = 32'h4cc48e82;
    ram_cell[    2379] = 32'h653c1165;
    ram_cell[    2380] = 32'h88d99b22;
    ram_cell[    2381] = 32'hb41c7a6a;
    ram_cell[    2382] = 32'h18e2c6ea;
    ram_cell[    2383] = 32'h88454bcb;
    ram_cell[    2384] = 32'h77200328;
    ram_cell[    2385] = 32'hf860a27a;
    ram_cell[    2386] = 32'h467e3d61;
    ram_cell[    2387] = 32'hd3faabbb;
    ram_cell[    2388] = 32'hc5db5a01;
    ram_cell[    2389] = 32'he27400f6;
    ram_cell[    2390] = 32'h5bd944ed;
    ram_cell[    2391] = 32'h5f771ebe;
    ram_cell[    2392] = 32'h0c73aead;
    ram_cell[    2393] = 32'h1c19389e;
    ram_cell[    2394] = 32'ha2a5f70f;
    ram_cell[    2395] = 32'hf663eb8d;
    ram_cell[    2396] = 32'ha39b62f6;
    ram_cell[    2397] = 32'h76afbcd2;
    ram_cell[    2398] = 32'h24db9ea4;
    ram_cell[    2399] = 32'hd7d39a87;
    ram_cell[    2400] = 32'h933241fd;
    ram_cell[    2401] = 32'h385738c5;
    ram_cell[    2402] = 32'h66682293;
    ram_cell[    2403] = 32'h21a5eb24;
    ram_cell[    2404] = 32'hf1e905bc;
    ram_cell[    2405] = 32'h5e0797f5;
    ram_cell[    2406] = 32'h2ad1d604;
    ram_cell[    2407] = 32'h1db391cd;
    ram_cell[    2408] = 32'h45fbe1c9;
    ram_cell[    2409] = 32'h93bbcbc2;
    ram_cell[    2410] = 32'h0ba8fe42;
    ram_cell[    2411] = 32'h4b9e4c33;
    ram_cell[    2412] = 32'haa3d6869;
    ram_cell[    2413] = 32'hf9426a03;
    ram_cell[    2414] = 32'h7da60694;
    ram_cell[    2415] = 32'hf4e5c7c0;
    ram_cell[    2416] = 32'hdc4128e1;
    ram_cell[    2417] = 32'h75307a02;
    ram_cell[    2418] = 32'hed00d20e;
    ram_cell[    2419] = 32'h9c30bf9d;
    ram_cell[    2420] = 32'h52a677f5;
    ram_cell[    2421] = 32'hbf52e4a9;
    ram_cell[    2422] = 32'h7c899390;
    ram_cell[    2423] = 32'h6f1af0c7;
    ram_cell[    2424] = 32'hdb4f72cb;
    ram_cell[    2425] = 32'h2cef37d2;
    ram_cell[    2426] = 32'h44e05904;
    ram_cell[    2427] = 32'hed81dcff;
    ram_cell[    2428] = 32'h015cfb35;
    ram_cell[    2429] = 32'hf279e52c;
    ram_cell[    2430] = 32'ha9fa2e00;
    ram_cell[    2431] = 32'hc383f5e1;
    ram_cell[    2432] = 32'h86c509dc;
    ram_cell[    2433] = 32'h470066fe;
    ram_cell[    2434] = 32'h2a531313;
    ram_cell[    2435] = 32'hf1c9060d;
    ram_cell[    2436] = 32'h3653157f;
    ram_cell[    2437] = 32'h529b5b77;
    ram_cell[    2438] = 32'hce14c91f;
    ram_cell[    2439] = 32'hb0187a99;
    ram_cell[    2440] = 32'hd123bc23;
    ram_cell[    2441] = 32'h6ad34b3a;
    ram_cell[    2442] = 32'h62b998ec;
    ram_cell[    2443] = 32'hd25cc9c3;
    ram_cell[    2444] = 32'ha3b7e639;
    ram_cell[    2445] = 32'hf4194ec6;
    ram_cell[    2446] = 32'h55c83fd1;
    ram_cell[    2447] = 32'hc92e0bff;
    ram_cell[    2448] = 32'hbf2062cd;
    ram_cell[    2449] = 32'hcc88077a;
    ram_cell[    2450] = 32'hb0211e32;
    ram_cell[    2451] = 32'h3e134d67;
    ram_cell[    2452] = 32'h9d2ff245;
    ram_cell[    2453] = 32'h6247565b;
    ram_cell[    2454] = 32'h1b0456e5;
    ram_cell[    2455] = 32'had9227f5;
    ram_cell[    2456] = 32'h9f60db45;
    ram_cell[    2457] = 32'h6aff8546;
    ram_cell[    2458] = 32'h93cbf633;
    ram_cell[    2459] = 32'hb3094f25;
    ram_cell[    2460] = 32'haeebdb48;
    ram_cell[    2461] = 32'h5f4badbc;
    ram_cell[    2462] = 32'h689dcc76;
    ram_cell[    2463] = 32'h80c6488d;
    ram_cell[    2464] = 32'h01276ed1;
    ram_cell[    2465] = 32'h3cb6897e;
    ram_cell[    2466] = 32'h83d5ffeb;
    ram_cell[    2467] = 32'h6b10931a;
    ram_cell[    2468] = 32'hc8d64f99;
    ram_cell[    2469] = 32'h8c48dbec;
    ram_cell[    2470] = 32'h2d99e02e;
    ram_cell[    2471] = 32'hbf18b25d;
    ram_cell[    2472] = 32'h9f46c634;
    ram_cell[    2473] = 32'h4384d676;
    ram_cell[    2474] = 32'hc20591d4;
    ram_cell[    2475] = 32'h1d913be6;
    ram_cell[    2476] = 32'h52ecba9e;
    ram_cell[    2477] = 32'ha0d269d8;
    ram_cell[    2478] = 32'h1568b164;
    ram_cell[    2479] = 32'h9fa87fda;
    ram_cell[    2480] = 32'hc92a0884;
    ram_cell[    2481] = 32'h30be6f2f;
    ram_cell[    2482] = 32'h5a313040;
    ram_cell[    2483] = 32'hb85b4ed3;
    ram_cell[    2484] = 32'h97d30365;
    ram_cell[    2485] = 32'h401e7332;
    ram_cell[    2486] = 32'h92afc104;
    ram_cell[    2487] = 32'hc05f51c4;
    ram_cell[    2488] = 32'h6cbf05b3;
    ram_cell[    2489] = 32'h5918f1fb;
    ram_cell[    2490] = 32'h3e23b93f;
    ram_cell[    2491] = 32'hd51b4ec0;
    ram_cell[    2492] = 32'h4f2ef860;
    ram_cell[    2493] = 32'h2baba16b;
    ram_cell[    2494] = 32'hb9ea1948;
    ram_cell[    2495] = 32'h3ead36c0;
    ram_cell[    2496] = 32'h75cefd52;
    ram_cell[    2497] = 32'h96d2582d;
    ram_cell[    2498] = 32'he414f47c;
    ram_cell[    2499] = 32'hd661e7cb;
    ram_cell[    2500] = 32'h4dd60031;
    ram_cell[    2501] = 32'h27b87cbe;
    ram_cell[    2502] = 32'he0124340;
    ram_cell[    2503] = 32'h0165029e;
    ram_cell[    2504] = 32'h1bbab8aa;
    ram_cell[    2505] = 32'hc29bc09b;
    ram_cell[    2506] = 32'h777cb2ea;
    ram_cell[    2507] = 32'h0249a42a;
    ram_cell[    2508] = 32'hb892a552;
    ram_cell[    2509] = 32'h2c6b5003;
    ram_cell[    2510] = 32'h9454f0d1;
    ram_cell[    2511] = 32'hb070a207;
    ram_cell[    2512] = 32'hebad2408;
    ram_cell[    2513] = 32'hef4761f3;
    ram_cell[    2514] = 32'he3ee29fc;
    ram_cell[    2515] = 32'hbb73856a;
    ram_cell[    2516] = 32'h8b16c51f;
    ram_cell[    2517] = 32'h33b1f8a2;
    ram_cell[    2518] = 32'h725292de;
    ram_cell[    2519] = 32'h7938e750;
    ram_cell[    2520] = 32'hcaf073f8;
    ram_cell[    2521] = 32'h9902e735;
    ram_cell[    2522] = 32'hd919e551;
    ram_cell[    2523] = 32'h9b951573;
    ram_cell[    2524] = 32'h87e6f9f2;
    ram_cell[    2525] = 32'h131bba44;
    ram_cell[    2526] = 32'heba77f3a;
    ram_cell[    2527] = 32'hefb77320;
    ram_cell[    2528] = 32'h5c43a6f9;
    ram_cell[    2529] = 32'h876cdc5d;
    ram_cell[    2530] = 32'h104552bc;
    ram_cell[    2531] = 32'ha7e9fa28;
    ram_cell[    2532] = 32'h8dc9b7d4;
    ram_cell[    2533] = 32'h6680e5c9;
    ram_cell[    2534] = 32'hb183dc0a;
    ram_cell[    2535] = 32'h3acd7f1a;
    ram_cell[    2536] = 32'hf2668c52;
    ram_cell[    2537] = 32'h467b79cb;
    ram_cell[    2538] = 32'h0df5d16e;
    ram_cell[    2539] = 32'h000fe728;
    ram_cell[    2540] = 32'hfd40b94a;
    ram_cell[    2541] = 32'h34893ab2;
    ram_cell[    2542] = 32'hdf0ac6f6;
    ram_cell[    2543] = 32'hd11e8eec;
    ram_cell[    2544] = 32'h45588b7d;
    ram_cell[    2545] = 32'ha9e44493;
    ram_cell[    2546] = 32'h7ed82e11;
    ram_cell[    2547] = 32'hacd14b89;
    ram_cell[    2548] = 32'h146ef3e4;
    ram_cell[    2549] = 32'hdea763c0;
    ram_cell[    2550] = 32'h8d02801c;
    ram_cell[    2551] = 32'hf7a598ef;
    ram_cell[    2552] = 32'h169209c8;
    ram_cell[    2553] = 32'hd372d97f;
    ram_cell[    2554] = 32'h78a4bc14;
    ram_cell[    2555] = 32'h3813fb11;
    ram_cell[    2556] = 32'h80ee89f3;
    ram_cell[    2557] = 32'h72e753b1;
    ram_cell[    2558] = 32'h20f652d4;
    ram_cell[    2559] = 32'h3356e3fe;
    ram_cell[    2560] = 32'h278440f1;
    ram_cell[    2561] = 32'h68a09cdf;
    ram_cell[    2562] = 32'h573f9a4c;
    ram_cell[    2563] = 32'h4e7f1527;
    ram_cell[    2564] = 32'h9c028dfa;
    ram_cell[    2565] = 32'ha79b3aa2;
    ram_cell[    2566] = 32'ha42c2670;
    ram_cell[    2567] = 32'he756e7b7;
    ram_cell[    2568] = 32'hcc668811;
    ram_cell[    2569] = 32'h4e1f9ef5;
    ram_cell[    2570] = 32'h17522828;
    ram_cell[    2571] = 32'hbf154bbd;
    ram_cell[    2572] = 32'hbe00f937;
    ram_cell[    2573] = 32'h44941579;
    ram_cell[    2574] = 32'h893c79a6;
    ram_cell[    2575] = 32'he54ff20b;
    ram_cell[    2576] = 32'ha4a4136e;
    ram_cell[    2577] = 32'h15d38c2d;
    ram_cell[    2578] = 32'h13928c2c;
    ram_cell[    2579] = 32'h3f7c47b6;
    ram_cell[    2580] = 32'hffa0969b;
    ram_cell[    2581] = 32'h225bca8e;
    ram_cell[    2582] = 32'h298c2440;
    ram_cell[    2583] = 32'h98ffc7ec;
    ram_cell[    2584] = 32'h038310ed;
    ram_cell[    2585] = 32'h80bae575;
    ram_cell[    2586] = 32'hd4ae2b92;
    ram_cell[    2587] = 32'h0192a19f;
    ram_cell[    2588] = 32'h581f6206;
    ram_cell[    2589] = 32'hc8f03272;
    ram_cell[    2590] = 32'ha67fc0ca;
    ram_cell[    2591] = 32'h741dbeb8;
    ram_cell[    2592] = 32'hc09c40a5;
    ram_cell[    2593] = 32'hb50aad45;
    ram_cell[    2594] = 32'h7d89411b;
    ram_cell[    2595] = 32'hc381cc73;
    ram_cell[    2596] = 32'h00d2e121;
    ram_cell[    2597] = 32'he8e5e140;
    ram_cell[    2598] = 32'hf1c49a79;
    ram_cell[    2599] = 32'h9f146091;
    ram_cell[    2600] = 32'h6aba733f;
    ram_cell[    2601] = 32'h91658df4;
    ram_cell[    2602] = 32'h8e2d715e;
    ram_cell[    2603] = 32'h1b1221b0;
    ram_cell[    2604] = 32'h4ec53e3e;
    ram_cell[    2605] = 32'h7e91573a;
    ram_cell[    2606] = 32'h2c755428;
    ram_cell[    2607] = 32'h9525b27b;
    ram_cell[    2608] = 32'h7cf00fec;
    ram_cell[    2609] = 32'h63739ada;
    ram_cell[    2610] = 32'hb23368d6;
    ram_cell[    2611] = 32'h510d1cad;
    ram_cell[    2612] = 32'h4651982a;
    ram_cell[    2613] = 32'h6a6b5c5a;
    ram_cell[    2614] = 32'h75d0be3e;
    ram_cell[    2615] = 32'haecfb5c1;
    ram_cell[    2616] = 32'h7849efb5;
    ram_cell[    2617] = 32'hae4d5195;
    ram_cell[    2618] = 32'hd4a33cbb;
    ram_cell[    2619] = 32'h6fe244f4;
    ram_cell[    2620] = 32'h29dc82b6;
    ram_cell[    2621] = 32'hc5e9fe4c;
    ram_cell[    2622] = 32'h1ff43366;
    ram_cell[    2623] = 32'h2cbed160;
    ram_cell[    2624] = 32'h9199888c;
    ram_cell[    2625] = 32'h99597015;
    ram_cell[    2626] = 32'h495c4e08;
    ram_cell[    2627] = 32'hfd0eb486;
    ram_cell[    2628] = 32'h580357a3;
    ram_cell[    2629] = 32'h74c30b89;
    ram_cell[    2630] = 32'h696d45b0;
    ram_cell[    2631] = 32'h8b379c3d;
    ram_cell[    2632] = 32'h271755e2;
    ram_cell[    2633] = 32'h156ba897;
    ram_cell[    2634] = 32'hef0c0fe5;
    ram_cell[    2635] = 32'hda63d209;
    ram_cell[    2636] = 32'h1d483bad;
    ram_cell[    2637] = 32'h57186ca9;
    ram_cell[    2638] = 32'hfad21b8e;
    ram_cell[    2639] = 32'hd18a5ab7;
    ram_cell[    2640] = 32'hd59a7964;
    ram_cell[    2641] = 32'h22461f80;
    ram_cell[    2642] = 32'hccc21d67;
    ram_cell[    2643] = 32'hb6abe28d;
    ram_cell[    2644] = 32'h32b184bb;
    ram_cell[    2645] = 32'hfea3f404;
    ram_cell[    2646] = 32'h35c627d9;
    ram_cell[    2647] = 32'h46bc3480;
    ram_cell[    2648] = 32'h6031b5c8;
    ram_cell[    2649] = 32'h2c1ea3b6;
    ram_cell[    2650] = 32'h1abafc54;
    ram_cell[    2651] = 32'hfcc45b54;
    ram_cell[    2652] = 32'h0a62cef6;
    ram_cell[    2653] = 32'h7c8c9171;
    ram_cell[    2654] = 32'ha378f8e8;
    ram_cell[    2655] = 32'h5f4c4ef7;
    ram_cell[    2656] = 32'h71bff2f6;
    ram_cell[    2657] = 32'h0f3ccd69;
    ram_cell[    2658] = 32'h08bd5bb7;
    ram_cell[    2659] = 32'h01b9fe06;
    ram_cell[    2660] = 32'hbbc7c5a4;
    ram_cell[    2661] = 32'hc5a38271;
    ram_cell[    2662] = 32'h556bb5f5;
    ram_cell[    2663] = 32'heba9ddc6;
    ram_cell[    2664] = 32'hb7792a96;
    ram_cell[    2665] = 32'h3d0f09f9;
    ram_cell[    2666] = 32'hbc31a7fc;
    ram_cell[    2667] = 32'hd93135c8;
    ram_cell[    2668] = 32'h249b29c3;
    ram_cell[    2669] = 32'h8c36d50c;
    ram_cell[    2670] = 32'h5f3c921d;
    ram_cell[    2671] = 32'he1782a64;
    ram_cell[    2672] = 32'h9a1dd45c;
    ram_cell[    2673] = 32'h5c338413;
    ram_cell[    2674] = 32'hee13d71c;
    ram_cell[    2675] = 32'hfe2eacd7;
    ram_cell[    2676] = 32'h3efddf34;
    ram_cell[    2677] = 32'h8f387e0d;
    ram_cell[    2678] = 32'h2e9c2ff8;
    ram_cell[    2679] = 32'h8bd2b549;
    ram_cell[    2680] = 32'h1a97eaf2;
    ram_cell[    2681] = 32'h3385344b;
    ram_cell[    2682] = 32'ha9d05f9f;
    ram_cell[    2683] = 32'hd16c9e23;
    ram_cell[    2684] = 32'h2262ee64;
    ram_cell[    2685] = 32'h06e6b02f;
    ram_cell[    2686] = 32'h8e3d9ad7;
    ram_cell[    2687] = 32'h853de827;
    ram_cell[    2688] = 32'hd9df4d6f;
    ram_cell[    2689] = 32'h5adc1bff;
    ram_cell[    2690] = 32'hab6a3709;
    ram_cell[    2691] = 32'h5dfa852b;
    ram_cell[    2692] = 32'hf5041012;
    ram_cell[    2693] = 32'h786cb61e;
    ram_cell[    2694] = 32'haf9aea60;
    ram_cell[    2695] = 32'h7e2eeb42;
    ram_cell[    2696] = 32'h4d1f2ac9;
    ram_cell[    2697] = 32'h42e6e3cc;
    ram_cell[    2698] = 32'h66f5f14d;
    ram_cell[    2699] = 32'h61bb552d;
    ram_cell[    2700] = 32'h1d2ab8cf;
    ram_cell[    2701] = 32'ha843db0d;
    ram_cell[    2702] = 32'hd3e8a3c5;
    ram_cell[    2703] = 32'h61036566;
    ram_cell[    2704] = 32'hccf477e1;
    ram_cell[    2705] = 32'hf9e66a2d;
    ram_cell[    2706] = 32'h8e874de8;
    ram_cell[    2707] = 32'h350400e8;
    ram_cell[    2708] = 32'h964bbb64;
    ram_cell[    2709] = 32'h0d532a1c;
    ram_cell[    2710] = 32'hc47d25a2;
    ram_cell[    2711] = 32'he28771b5;
    ram_cell[    2712] = 32'hb940a0a3;
    ram_cell[    2713] = 32'he3424c96;
    ram_cell[    2714] = 32'h6939bf70;
    ram_cell[    2715] = 32'h991fcfbb;
    ram_cell[    2716] = 32'h537b93bf;
    ram_cell[    2717] = 32'ha7dac465;
    ram_cell[    2718] = 32'h068f1127;
    ram_cell[    2719] = 32'h024f3c92;
    ram_cell[    2720] = 32'hebe925e9;
    ram_cell[    2721] = 32'h2f36db15;
    ram_cell[    2722] = 32'h0da3b2e0;
    ram_cell[    2723] = 32'h8910dae3;
    ram_cell[    2724] = 32'h59a5458d;
    ram_cell[    2725] = 32'ha13e13f3;
    ram_cell[    2726] = 32'h01c89cd7;
    ram_cell[    2727] = 32'hc1caab96;
    ram_cell[    2728] = 32'h57b435f8;
    ram_cell[    2729] = 32'h1b812a2f;
    ram_cell[    2730] = 32'h4cd588ee;
    ram_cell[    2731] = 32'h8fa7cc72;
    ram_cell[    2732] = 32'hee5ab673;
    ram_cell[    2733] = 32'h81bb6437;
    ram_cell[    2734] = 32'h45f0cdef;
    ram_cell[    2735] = 32'hea4603f9;
    ram_cell[    2736] = 32'hefbeaf11;
    ram_cell[    2737] = 32'h9852143b;
    ram_cell[    2738] = 32'hb2c293f8;
    ram_cell[    2739] = 32'he8d70d7c;
    ram_cell[    2740] = 32'h08562288;
    ram_cell[    2741] = 32'h286fb17f;
    ram_cell[    2742] = 32'hb8880fec;
    ram_cell[    2743] = 32'he89f0083;
    ram_cell[    2744] = 32'h24a2e32d;
    ram_cell[    2745] = 32'h03c2f77b;
    ram_cell[    2746] = 32'h2d5b6a4d;
    ram_cell[    2747] = 32'he4405ffd;
    ram_cell[    2748] = 32'hf725415d;
    ram_cell[    2749] = 32'h94c73f15;
    ram_cell[    2750] = 32'h5c14146c;
    ram_cell[    2751] = 32'h084a26a6;
    ram_cell[    2752] = 32'h7a35f781;
    ram_cell[    2753] = 32'h034fa2b9;
    ram_cell[    2754] = 32'h17e50676;
    ram_cell[    2755] = 32'h8a697b1f;
    ram_cell[    2756] = 32'hdc4386f0;
    ram_cell[    2757] = 32'h08adf7ed;
    ram_cell[    2758] = 32'h67195c24;
    ram_cell[    2759] = 32'h9adc5fcc;
    ram_cell[    2760] = 32'h093c18cb;
    ram_cell[    2761] = 32'hefeaa7e3;
    ram_cell[    2762] = 32'h8275c8ef;
    ram_cell[    2763] = 32'h1f3cf3de;
    ram_cell[    2764] = 32'h149d304a;
    ram_cell[    2765] = 32'h4e3e626b;
    ram_cell[    2766] = 32'h0e300446;
    ram_cell[    2767] = 32'hd1de4992;
    ram_cell[    2768] = 32'h69c533ac;
    ram_cell[    2769] = 32'h6ab2e4ce;
    ram_cell[    2770] = 32'hc249eda2;
    ram_cell[    2771] = 32'hb24ad6c9;
    ram_cell[    2772] = 32'he2014681;
    ram_cell[    2773] = 32'hcf3334ae;
    ram_cell[    2774] = 32'h93e84843;
    ram_cell[    2775] = 32'h2f9e9a9b;
    ram_cell[    2776] = 32'h8a827fd5;
    ram_cell[    2777] = 32'hf4cdb1e6;
    ram_cell[    2778] = 32'h43d93f35;
    ram_cell[    2779] = 32'h8de15bfa;
    ram_cell[    2780] = 32'h2cb9396f;
    ram_cell[    2781] = 32'hc3889fa7;
    ram_cell[    2782] = 32'h20380cfe;
    ram_cell[    2783] = 32'h692e5179;
    ram_cell[    2784] = 32'h1a0571b4;
    ram_cell[    2785] = 32'hfea11006;
    ram_cell[    2786] = 32'h01e7e41b;
    ram_cell[    2787] = 32'h4201fdb5;
    ram_cell[    2788] = 32'hdd590e39;
    ram_cell[    2789] = 32'h03d2078d;
    ram_cell[    2790] = 32'h00301877;
    ram_cell[    2791] = 32'h1d09afc2;
    ram_cell[    2792] = 32'hf662207a;
    ram_cell[    2793] = 32'hcfc63a8a;
    ram_cell[    2794] = 32'h316694e7;
    ram_cell[    2795] = 32'hffeadeb2;
    ram_cell[    2796] = 32'h2f0a836b;
    ram_cell[    2797] = 32'h0e7a54fb;
    ram_cell[    2798] = 32'h20c9580d;
    ram_cell[    2799] = 32'h34a469f5;
    ram_cell[    2800] = 32'hd0cdad9d;
    ram_cell[    2801] = 32'hfb8ba122;
    ram_cell[    2802] = 32'h5486c708;
    ram_cell[    2803] = 32'hd5782b5d;
    ram_cell[    2804] = 32'h0642ae66;
    ram_cell[    2805] = 32'hcfbd3ae0;
    ram_cell[    2806] = 32'h08cebda8;
    ram_cell[    2807] = 32'hd64624f7;
    ram_cell[    2808] = 32'h274a8ab9;
    ram_cell[    2809] = 32'hf99e0bda;
    ram_cell[    2810] = 32'h50f23a05;
    ram_cell[    2811] = 32'ha82fc3a5;
    ram_cell[    2812] = 32'he70fe100;
    ram_cell[    2813] = 32'h5ea0dc87;
    ram_cell[    2814] = 32'h201ab68c;
    ram_cell[    2815] = 32'h58b36885;
    ram_cell[    2816] = 32'h673c5056;
    ram_cell[    2817] = 32'h42576075;
    ram_cell[    2818] = 32'h36fe04e7;
    ram_cell[    2819] = 32'ha300310d;
    ram_cell[    2820] = 32'hec8e2b54;
    ram_cell[    2821] = 32'h832c6fe6;
    ram_cell[    2822] = 32'h86e5c11c;
    ram_cell[    2823] = 32'he8cbdbb2;
    ram_cell[    2824] = 32'h57f9e4b7;
    ram_cell[    2825] = 32'h26b0b482;
    ram_cell[    2826] = 32'h63914ba8;
    ram_cell[    2827] = 32'h28770669;
    ram_cell[    2828] = 32'h70c377ab;
    ram_cell[    2829] = 32'hb513abf9;
    ram_cell[    2830] = 32'h20b22549;
    ram_cell[    2831] = 32'h572f1bc3;
    ram_cell[    2832] = 32'h8c2d38bc;
    ram_cell[    2833] = 32'h3eda6dac;
    ram_cell[    2834] = 32'hf0559171;
    ram_cell[    2835] = 32'h0ce61a8c;
    ram_cell[    2836] = 32'h9dd20891;
    ram_cell[    2837] = 32'hf988f676;
    ram_cell[    2838] = 32'h89795aad;
    ram_cell[    2839] = 32'h9ebc8e06;
    ram_cell[    2840] = 32'h9534459c;
    ram_cell[    2841] = 32'ha35cc985;
    ram_cell[    2842] = 32'h65de62cd;
    ram_cell[    2843] = 32'hc6471e08;
    ram_cell[    2844] = 32'h34ca2f03;
    ram_cell[    2845] = 32'h408cf749;
    ram_cell[    2846] = 32'hb3ac5f77;
    ram_cell[    2847] = 32'ha83e8aca;
    ram_cell[    2848] = 32'he97e6227;
    ram_cell[    2849] = 32'h2bb6847d;
    ram_cell[    2850] = 32'h04d53502;
    ram_cell[    2851] = 32'h69db90f6;
    ram_cell[    2852] = 32'h593ae0f9;
    ram_cell[    2853] = 32'hba7a37c0;
    ram_cell[    2854] = 32'h7dced4e0;
    ram_cell[    2855] = 32'ha46b413c;
    ram_cell[    2856] = 32'hb7c61ec5;
    ram_cell[    2857] = 32'h39d28f44;
    ram_cell[    2858] = 32'h3c3c0c94;
    ram_cell[    2859] = 32'h94d5f835;
    ram_cell[    2860] = 32'hda45f2be;
    ram_cell[    2861] = 32'h5491b034;
    ram_cell[    2862] = 32'h2fe24140;
    ram_cell[    2863] = 32'hadb21059;
    ram_cell[    2864] = 32'hd3ad3636;
    ram_cell[    2865] = 32'hb86f521c;
    ram_cell[    2866] = 32'h26533373;
    ram_cell[    2867] = 32'h1f07c6bf;
    ram_cell[    2868] = 32'h83f82e29;
    ram_cell[    2869] = 32'he6e95aac;
    ram_cell[    2870] = 32'h31589049;
    ram_cell[    2871] = 32'hb9d7ffb1;
    ram_cell[    2872] = 32'h7de9ca46;
    ram_cell[    2873] = 32'h859164d7;
    ram_cell[    2874] = 32'hcbaf378f;
    ram_cell[    2875] = 32'h371ec0b0;
    ram_cell[    2876] = 32'ha5da25b2;
    ram_cell[    2877] = 32'h9552985e;
    ram_cell[    2878] = 32'h69615462;
    ram_cell[    2879] = 32'h3800816e;
    ram_cell[    2880] = 32'h137dd962;
    ram_cell[    2881] = 32'h641052de;
    ram_cell[    2882] = 32'h44c65df8;
    ram_cell[    2883] = 32'hc2e4cf1f;
    ram_cell[    2884] = 32'h9ec6dbfb;
    ram_cell[    2885] = 32'hdd1f797b;
    ram_cell[    2886] = 32'hebaf438f;
    ram_cell[    2887] = 32'hbcae6bc2;
    ram_cell[    2888] = 32'h155769ba;
    ram_cell[    2889] = 32'h99de577c;
    ram_cell[    2890] = 32'hfce13b3f;
    ram_cell[    2891] = 32'h7494cfae;
    ram_cell[    2892] = 32'h2e8b3c93;
    ram_cell[    2893] = 32'h5229450d;
    ram_cell[    2894] = 32'h52e62708;
    ram_cell[    2895] = 32'hb110b146;
    ram_cell[    2896] = 32'h271117f1;
    ram_cell[    2897] = 32'h06117917;
    ram_cell[    2898] = 32'h3ac0a05d;
    ram_cell[    2899] = 32'h3dfe2248;
    ram_cell[    2900] = 32'hd9c2a539;
    ram_cell[    2901] = 32'h2d11e91c;
    ram_cell[    2902] = 32'h5e0ccf59;
    ram_cell[    2903] = 32'h5ca8f23f;
    ram_cell[    2904] = 32'h9e9abcf6;
    ram_cell[    2905] = 32'hd4b3279c;
    ram_cell[    2906] = 32'h99c117c1;
    ram_cell[    2907] = 32'h81de8431;
    ram_cell[    2908] = 32'hcb7c66d0;
    ram_cell[    2909] = 32'h529f03cc;
    ram_cell[    2910] = 32'haac75b75;
    ram_cell[    2911] = 32'h664c4623;
    ram_cell[    2912] = 32'hd4cfac73;
    ram_cell[    2913] = 32'h273eca7f;
    ram_cell[    2914] = 32'h881bcb8a;
    ram_cell[    2915] = 32'h65fde6b0;
    ram_cell[    2916] = 32'he7d9e251;
    ram_cell[    2917] = 32'h0e70b4af;
    ram_cell[    2918] = 32'h5571827b;
    ram_cell[    2919] = 32'h967f5472;
    ram_cell[    2920] = 32'hf5a3bcec;
    ram_cell[    2921] = 32'h9100df41;
    ram_cell[    2922] = 32'h0f43c74f;
    ram_cell[    2923] = 32'h6fcac071;
    ram_cell[    2924] = 32'h9474481b;
    ram_cell[    2925] = 32'heb1c637e;
    ram_cell[    2926] = 32'h8825dd7e;
    ram_cell[    2927] = 32'h957fd785;
    ram_cell[    2928] = 32'ha902475f;
    ram_cell[    2929] = 32'h5f3c9993;
    ram_cell[    2930] = 32'hfa7b30c1;
    ram_cell[    2931] = 32'h97682eb9;
    ram_cell[    2932] = 32'hf95016db;
    ram_cell[    2933] = 32'h0ef6b070;
    ram_cell[    2934] = 32'h66337bd0;
    ram_cell[    2935] = 32'h89928553;
    ram_cell[    2936] = 32'h9630eacd;
    ram_cell[    2937] = 32'h3e827ddd;
    ram_cell[    2938] = 32'h23439ace;
    ram_cell[    2939] = 32'hf712f4cb;
    ram_cell[    2940] = 32'hac8181b8;
    ram_cell[    2941] = 32'h04c99bb6;
    ram_cell[    2942] = 32'hcf6a5d7a;
    ram_cell[    2943] = 32'hda41d4e8;
    ram_cell[    2944] = 32'hb6d17992;
    ram_cell[    2945] = 32'h031145e5;
    ram_cell[    2946] = 32'h30ae0e60;
    ram_cell[    2947] = 32'he20739b9;
    ram_cell[    2948] = 32'h64b12817;
    ram_cell[    2949] = 32'h2f200dc1;
    ram_cell[    2950] = 32'h4d40c688;
    ram_cell[    2951] = 32'h96086e47;
    ram_cell[    2952] = 32'h6f974645;
    ram_cell[    2953] = 32'h476e25b3;
    ram_cell[    2954] = 32'h6e24626c;
    ram_cell[    2955] = 32'h8be42bd3;
    ram_cell[    2956] = 32'hdd85c4a3;
    ram_cell[    2957] = 32'he10784b0;
    ram_cell[    2958] = 32'h4237dab4;
    ram_cell[    2959] = 32'h8a23cbb9;
    ram_cell[    2960] = 32'hfb42814d;
    ram_cell[    2961] = 32'h99ee7077;
    ram_cell[    2962] = 32'h47cf2866;
    ram_cell[    2963] = 32'hdb394745;
    ram_cell[    2964] = 32'h78ec7bd0;
    ram_cell[    2965] = 32'hd219edd4;
    ram_cell[    2966] = 32'hdbb3abb3;
    ram_cell[    2967] = 32'h188ce02e;
    ram_cell[    2968] = 32'ha5e88856;
    ram_cell[    2969] = 32'ha70f4879;
    ram_cell[    2970] = 32'h95e6086b;
    ram_cell[    2971] = 32'hbae7240b;
    ram_cell[    2972] = 32'h26aa12f4;
    ram_cell[    2973] = 32'h4d2c1869;
    ram_cell[    2974] = 32'h7f6a1338;
    ram_cell[    2975] = 32'h6b146ce5;
    ram_cell[    2976] = 32'h1b6e05ba;
    ram_cell[    2977] = 32'hfdb6eae3;
    ram_cell[    2978] = 32'ha74ced5d;
    ram_cell[    2979] = 32'hfc31910d;
    ram_cell[    2980] = 32'hdf45ee94;
    ram_cell[    2981] = 32'hf0d9d1a4;
    ram_cell[    2982] = 32'h006f6bb9;
    ram_cell[    2983] = 32'h343e8515;
    ram_cell[    2984] = 32'h154a4b98;
    ram_cell[    2985] = 32'h5855d33c;
    ram_cell[    2986] = 32'hec04090c;
    ram_cell[    2987] = 32'h13c3fa1b;
    ram_cell[    2988] = 32'h4c3dcd97;
    ram_cell[    2989] = 32'haca9dbfa;
    ram_cell[    2990] = 32'hb7b45b4a;
    ram_cell[    2991] = 32'h312c460f;
    ram_cell[    2992] = 32'ha34e13f3;
    ram_cell[    2993] = 32'h5fc798bf;
    ram_cell[    2994] = 32'hc3e4afd2;
    ram_cell[    2995] = 32'hd47f2e29;
    ram_cell[    2996] = 32'h04ca7fbe;
    ram_cell[    2997] = 32'hefe52ff7;
    ram_cell[    2998] = 32'h052b862c;
    ram_cell[    2999] = 32'hda4899f4;
    ram_cell[    3000] = 32'h828b5940;
    ram_cell[    3001] = 32'hb94cdb8d;
    ram_cell[    3002] = 32'h99954144;
    ram_cell[    3003] = 32'h11254680;
    ram_cell[    3004] = 32'hffc03db8;
    ram_cell[    3005] = 32'h6193f915;
    ram_cell[    3006] = 32'hb443b091;
    ram_cell[    3007] = 32'h7d6a2b9b;
    ram_cell[    3008] = 32'ha996e733;
    ram_cell[    3009] = 32'hcde759ee;
    ram_cell[    3010] = 32'hf983a4e2;
    ram_cell[    3011] = 32'h9d6922ae;
    ram_cell[    3012] = 32'h5f807283;
    ram_cell[    3013] = 32'h628324b3;
    ram_cell[    3014] = 32'hb37d841c;
    ram_cell[    3015] = 32'h6e429c21;
    ram_cell[    3016] = 32'hfe7d8a47;
    ram_cell[    3017] = 32'h17454280;
    ram_cell[    3018] = 32'h1b842169;
    ram_cell[    3019] = 32'h6fe3007a;
    ram_cell[    3020] = 32'h59809fba;
    ram_cell[    3021] = 32'h9e302950;
    ram_cell[    3022] = 32'h3d35689d;
    ram_cell[    3023] = 32'h6579380a;
    ram_cell[    3024] = 32'hc10fda7f;
    ram_cell[    3025] = 32'hfb15490b;
    ram_cell[    3026] = 32'he2cfde81;
    ram_cell[    3027] = 32'hbfcce9bb;
    ram_cell[    3028] = 32'hd9fd6ef9;
    ram_cell[    3029] = 32'hebf70c28;
    ram_cell[    3030] = 32'he6d4b3db;
    ram_cell[    3031] = 32'hb194c26a;
    ram_cell[    3032] = 32'hdf69e5ce;
    ram_cell[    3033] = 32'he2dc1764;
    ram_cell[    3034] = 32'ha5da08e0;
    ram_cell[    3035] = 32'h12390439;
    ram_cell[    3036] = 32'hfdf7b7ce;
    ram_cell[    3037] = 32'h874019fb;
    ram_cell[    3038] = 32'hfee72d17;
    ram_cell[    3039] = 32'ha59a102d;
    ram_cell[    3040] = 32'h4f02e77b;
    ram_cell[    3041] = 32'h8d8c2d96;
    ram_cell[    3042] = 32'h3020e8f8;
    ram_cell[    3043] = 32'hf0f8df88;
    ram_cell[    3044] = 32'h05cc6b4b;
    ram_cell[    3045] = 32'h4eee8d0e;
    ram_cell[    3046] = 32'hb27e7c7e;
    ram_cell[    3047] = 32'h62cac2e7;
    ram_cell[    3048] = 32'hccb966fe;
    ram_cell[    3049] = 32'he68ed362;
    ram_cell[    3050] = 32'h94729c96;
    ram_cell[    3051] = 32'h1219071a;
    ram_cell[    3052] = 32'h436be9b1;
    ram_cell[    3053] = 32'h21bf156e;
    ram_cell[    3054] = 32'h075314a9;
    ram_cell[    3055] = 32'h1049e129;
    ram_cell[    3056] = 32'h2cf6b7da;
    ram_cell[    3057] = 32'h5f21bd22;
    ram_cell[    3058] = 32'h194b672d;
    ram_cell[    3059] = 32'hd2f9dd28;
    ram_cell[    3060] = 32'h5ed25c82;
    ram_cell[    3061] = 32'h3eb61632;
    ram_cell[    3062] = 32'hd5ab1d23;
    ram_cell[    3063] = 32'h5021efc1;
    ram_cell[    3064] = 32'hda1c2934;
    ram_cell[    3065] = 32'h77789380;
    ram_cell[    3066] = 32'hd8e6278c;
    ram_cell[    3067] = 32'h4b9cb4e1;
    ram_cell[    3068] = 32'h9e773890;
    ram_cell[    3069] = 32'hdf4b9a1c;
    ram_cell[    3070] = 32'ha7e3641a;
    ram_cell[    3071] = 32'h7e1ad4be;
end

endmodule

